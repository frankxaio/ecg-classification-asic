module linear_tb;

    parameter MATRIX_SIZE = 16;
    parameter DATA_SIZE = 8;

    logic clk;
    logic reset;
    logic start;
    logic done;
    logic [DATA_SIZE-1:0] mat_a[MATRIX_SIZE-1:0][MATRIX_SIZE-1:0];
    logic [DATA_SIZE-1:0] wt[MATRIX_SIZE-1:0][MATRIX_SIZE-1:0];
    logic [DATA_SIZE-1:0] bias[MATRIX_SIZE-1:0];
    logic [DATA_SIZE-1:0] out_matrix[MATRIX_SIZE-1:0][MATRIX_SIZE-1:0];

    // 實例化linear模組
    linear #(
        .MATRIX_SIZE(MATRIX_SIZE),
        .DATA_SIZE  (DATA_SIZE)
    ) dut (
        .clk(clk),
        .reset(reset),
        .start(start),
        .done(done),
        .mat_a(mat_a),
        .wt(wt),
        .bias(bias),
        .out_matrix(out_matrix)
    );

    // 時脈生成
    always begin
        clk = 1'b0;
        #5;
        clk = 1'b1;
        #5;
    end

    // 測試激勵
    initial begin
        reset = 1'b1;
        start = 1'b0;
        #10;
        reset = 1'b0;
        #10;

        // 設定輸入矩陣和權重矩陣

        mat_a = '{
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1}
        };

        wt = '{
            '{2, 1, 3, 2, 1, 3, 2, 1, 3, 2, 1, 3, 2, 1, 3, 2},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{1, 3, 2, 1, 3, 2, 1, 3, 2, 1, 3, 2, 1, 3, 2, 1},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3},
            '{1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2},
            '{2, 1, 3, 2, 1, 3, 2, 1, 3, 2, 1, 3, 2, 1, 3, 2},
            '{2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2, 3, 1, 2}
        };

        bias = '{3, 1, 4, 2, 3, 1, 4, 2, 3, 1, 4, 2, 3, 1, 4, 2};

        #10;
        start = 1'b1;
        #10;
        start = 1'b0;

        wait (done);
        #10;

        // 檢查輸出矩陣
        for (int i = 0; i < MATRIX_SIZE; i++) begin
            for (int j = 0; j < MATRIX_SIZE; j++) begin
                $display("out_matrix[%0d][%0d] = %0d", i, j, out_matrix[i][j]);
            end
        end

        $finish;
    end

endmodule
