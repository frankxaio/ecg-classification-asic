module lut_module #(
    parameter ADDR_WIDTH = 8,
    parameter DATA_WIDTH = 8,
    parameter DATA_LEN   = 256
) (
    // input                                clk,
    // input                                rst,
    input               [ADDR_WIDTH-1:0] addr,
    output logic signed [DATA_WIDTH-1:0] data_o[0:DATA_LEN-1]
);


    localparam CLASSIFIER_BS_CNT = 6;
    localparam CLASSIFIER_WT_CNT = 96;
    localparam EMBEDDING_BS_CNT = 16;
    localparam EMBEDDING_WT_CNT = 16;
    localparam CLS_TOKEN_WT_CNT = 16;
    localparam FINAL_BS_CNT = 16;
    localparam FINAL_WT_CNT = 256;
    localparam KEYS_BS_CNT = 16;
    localparam KEYS_WT_CNT = 256;
    localparam QUERIES_BS_CNT = 16;
    localparam QUERIES_WT_CNT = 256;
    localparam VALUES_BS_CNT = 16;
    localparam VALUES_WT_CNT = 256;
    localparam MLP0_BS_CNT = 16;
    localparam MLP0_WT_CNT = 256;
    localparam MLP1_BS_CNT = 16;
    localparam MLP1_WT_CNT = 256;
    localparam PS_WT_CNT = 256;

    // Define the memory arrays for each file
    logic signed [DATA_WIDTH-1:0] classifier_bs[0:CLASSIFIER_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] classifier_wt[0:CLASSIFIER_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] embedding_bs[0:EMBEDDING_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] embedding_wt[0:EMBEDDING_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] cls_token_wt[0:CLS_TOKEN_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] final_bs[0:FINAL_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] final_wt[0:FINAL_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] keys_bs[0:KEYS_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] keys_wt[0:KEYS_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] queries_bs[0:QUERIES_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] queries_wt[0:QUERIES_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] values_bs[0:VALUES_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] values_wt[0:VALUES_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] mlp0_bs[0:MLP0_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] mlp0_wt[0:MLP0_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] mlp1_bs[0:MLP1_BS_CNT-1];
    logic signed [DATA_WIDTH-1:0] mlp1_wt[0:MLP1_WT_CNT-1];
    logic signed [DATA_WIDTH-1:0] ps_wt[0:PS_WT_CNT-1];

    // Array index register
    logic [$clog2(256):0] array_index, array_index_ns;
    logic [DATA_WIDTH-1:0] data;


    //LUT DATA
    assign classifier_bs = '{
            8'b00000100,
            8'b11111111,
            8'b00000000,
            8'b11111001,
            8'b00000000,
            8'b11111010
        };
    assign classifier_wt = '{
            8'b00000100,
            8'b11111011,
            8'b11111001,
            8'b11111010,
            8'b00000011,
            8'b11111000,
            8'b00001000,
            8'b00000111,
            8'b00000110,
            8'b00001000,
            8'b11111010,
            8'b00000000,
            8'b11111001,
            8'b00001000,
            8'b00000001,
            8'b00000000,
            8'b00001001,
            8'b00010010,
            8'b00001110,
            8'b11110101,
            8'b00001100,
            8'b00000100,
            8'b11101100,
            8'b00000010,
            8'b00000000,
            8'b00000011,
            8'b11110111,
            8'b00010110,
            8'b11111100,
            8'b11111111,
            8'b00001111,
            8'b11101101,
            8'b00001010,
            8'b11101101,
            8'b11111111,
            8'b00001110,
            8'b00000001,
            8'b00000001,
            8'b11111011,
            8'b11111011,
            8'b11110101,
            8'b11111010,
            8'b00001010,
            8'b00001110,
            8'b00000111,
            8'b11111000,
            8'b11111001,
            8'b00001011,
            8'b11111111,
            8'b11011000,
            8'b00001101,
            8'b00001101,
            8'b00001110,
            8'b00000100,
            8'b00000010,
            8'b11111110,
            8'b11111110,
            8'b11111010,
            8'b00000001,
            8'b11111101,
            8'b11111001,
            8'b00000010,
            8'b00000100,
            8'b00000010,
            8'b11110110,
            8'b00010010,
            8'b11101111,
            8'b00010100,
            8'b11101111,
            8'b00001111,
            8'b00000111,
            8'b11110011,
            8'b11110110,
            8'b11111001,
            8'b00001101,
            8'b11110001,
            8'b00001100,
            8'b11110001,
            8'b11110010,
            8'b11111010,
            8'b11111100,
            8'b00000111,
            8'b00001111,
            8'b11110110,
            8'b00000101,
            8'b00000110,
            8'b11111011,
            8'b00000110,
            8'b00000110,
            8'b00000011,
            8'b00000010,
            8'b11101101,
            8'b11111001,
            8'b00000011,
            8'b00000000,
            8'b00000101
        };
    assign embedding_bs = '{
            8'b11111010,
            8'b00010000,
            8'b11110010,
            8'b00001011,
            8'b11111101,
            8'b00000010,
            8'b11110101,
            8'b00001111,
            8'b00010001,
            8'b11111010,
            8'b00000000,
            8'b11110001,
            8'b00000111,
            8'b00001010,
            8'b00010001,
            8'b00000100
        };
    assign embedding_wt = '{
            8'b00001100,
            8'b11110001,
            8'b00001101,
            8'b11100100,
            8'b00000001,
            8'b00000101,
            8'b00000100,
            8'b00010110,
            8'b11101110,
            8'b11111101,
            8'b11111010,
            8'b11111101,
            8'b00010011,
            8'b11101000,
            8'b11011111,
            8'b00011011
        };
    assign cls_token_wt = '{
            8'b00000111,
            8'b00001111,
            8'b00000101,
            8'b11101001,
            8'b00001101,
            8'b00000100,
            8'b11111110,
            8'b00000011,
            8'b11111111,
            8'b11101101,
            8'b00010100,
            8'b00000011,
            8'b00000001,
            8'b00000110,
            8'b00001100,
            8'b00000110
        };
    assign final_bs = '{
            8'b00000011,
            8'b00000011,
            8'b11111100,
            8'b11111110,
            8'b11111101,
            8'b00000000,
            8'b11111110,
            8'b00000010,
            8'b00000110,
            8'b00000100,
            8'b00000010,
            8'b00000010,
            8'b11111111,
            8'b00000101,
            8'b00000010,
            8'b00000000
        };
    assign final_wt = '{
            8'b11111110,
            8'b00000010,
            8'b00000011,
            8'b00000110,
            8'b00000100,
            8'b00000111,
            8'b11111111,
            8'b11111111,
            8'b00000000,
            8'b00000100,
            8'b00000110,
            8'b11111111,
            8'b11111100,
            8'b00000100,
            8'b11111011,
            8'b00000101,
            8'b00000100,
            8'b00000000,
            8'b11111111,
            8'b00000111,
            8'b00000000,
            8'b11111101,
            8'b11111001,
            8'b00000101,
            8'b11111111,
            8'b11111011,
            8'b11111110,
            8'b00001000,
            8'b00000001,
            8'b00000011,
            8'b11111100,
            8'b00000000,
            8'b11111101,
            8'b11111110,
            8'b00000000,
            8'b00000011,
            8'b11111101,
            8'b00000010,
            8'b00000001,
            8'b11111101,
            8'b11111111,
            8'b00001110,
            8'b00000000,
            8'b11111101,
            8'b11111110,
            8'b00000100,
            8'b00000010,
            8'b00000001,
            8'b11111011,
            8'b11111110,
            8'b11111101,
            8'b11111101,
            8'b00000011,
            8'b00000000,
            8'b11111111,
            8'b00000000,
            8'b11111110,
            8'b00000011,
            8'b11111111,
            8'b11111111,
            8'b00000001,
            8'b00000010,
            8'b00000100,
            8'b00000101,
            8'b00000011,
            8'b00000011,
            8'b00000010,
            8'b11110111,
            8'b11111001,
            8'b00000010,
            8'b11111100,
            8'b11111011,
            8'b11111111,
            8'b00000111,
            8'b00000011,
            8'b11111100,
            8'b00000010,
            8'b11111100,
            8'b00000101,
            8'b00001110,
            8'b00000101,
            8'b00000000,
            8'b00000001,
            8'b11111100,
            8'b11101111,
            8'b00010111,
            8'b11101111,
            8'b11111101,
            8'b00000101,
            8'b00000100,
            8'b00000010,
            8'b00010001,
            8'b11111101,
            8'b00000100,
            8'b11111111,
            8'b00001010,
            8'b11111001,
            8'b00000011,
            8'b00000000,
            8'b00000011,
            8'b00000110,
            8'b00000001,
            8'b00000000,
            8'b11111100,
            8'b11111100,
            8'b00000001,
            8'b00000001,
            8'b00001001,
            8'b00000001,
            8'b11111011,
            8'b00000111,
            8'b11111011,
            8'b11111100,
            8'b00000100,
            8'b00000101,
            8'b00000101,
            8'b00000000,
            8'b00000001,
            8'b00000001,
            8'b11111110,
            8'b00000011,
            8'b00000000,
            8'b00000010,
            8'b00000010,
            8'b00000001,
            8'b00000001,
            8'b11111101,
            8'b11111011,
            8'b00000001,
            8'b00000101,
            8'b00001101,
            8'b00000100,
            8'b00000111,
            8'b00000101,
            8'b00001001,
            8'b11110110,
            8'b11111100,
            8'b00000111,
            8'b00001111,
            8'b00010100,
            8'b11110100,
            8'b11111011,
            8'b11111010,
            8'b11111001,
            8'b00000001,
            8'b00000111,
            8'b00000110,
            8'b00000001,
            8'b00000111,
            8'b00000101,
            8'b11111110,
            8'b00000000,
            8'b11111010,
            8'b00000110,
            8'b00000100,
            8'b00000000,
            8'b11111011,
            8'b00000001,
            8'b00000011,
            8'b00001000,
            8'b00000011,
            8'b11111100,
            8'b11111011,
            8'b11111000,
            8'b00000001,
            8'b00000111,
            8'b00000101,
            8'b00000101,
            8'b00000000,
            8'b00001001,
            8'b00000001,
            8'b11111100,
            8'b00000101,
            8'b00000011,
            8'b11111110,
            8'b00000000,
            8'b00000100,
            8'b00000010,
            8'b11111100,
            8'b11111101,
            8'b00000101,
            8'b11111011,
            8'b00000000,
            8'b00000001,
            8'b11111011,
            8'b11111011,
            8'b11111100,
            8'b11110001,
            8'b00000101,
            8'b11111101,
            8'b00000000,
            8'b00000101,
            8'b11111111,
            8'b11110111,
            8'b11101110,
            8'b11110111,
            8'b11111111,
            8'b00000101,
            8'b11110110,
            8'b00010101,
            8'b00001011,
            8'b00001010,
            8'b11110010,
            8'b11111001,
            8'b00001101,
            8'b00001100,
            8'b00000010,
            8'b00000111,
            8'b11111111,
            8'b00000101,
            8'b00001110,
            8'b00000100,
            8'b00000101,
            8'b11111101,
            8'b00001001,
            8'b11110110,
            8'b11110010,
            8'b00000001,
            8'b00001100,
            8'b00001000,
            8'b11110011,
            8'b11111000,
            8'b11111111,
            8'b11110100,
            8'b11111111,
            8'b00000101,
            8'b00001111,
            8'b00000110,
            8'b11111111,
            8'b11111110,
            8'b00000101,
            8'b11110100,
            8'b11111010,
            8'b11111111,
            8'b00001000,
            8'b00000100,
            8'b11111001,
            8'b11111001,
            8'b11111110,
            8'b00000001,
            8'b11111110,
            8'b00000001,
            8'b00000011,
            8'b00000011,
            8'b11111101,
            8'b11111111,
            8'b11111100,
            8'b11111110,
            8'b00000001,
            8'b11111000,
            8'b11111101,
            8'b00000000,
            8'b00000010,
            8'b11111110,
            8'b00000010,
            8'b00000101
        };
    assign keys_bs = '{
            8'b00000100,
            8'b11110111,
            8'b11111111,
            8'b11110011,
            8'b00000001,
            8'b11111111,
            8'b00000001,
            8'b00000001,
            8'b11111100,
            8'b00001001,
            8'b00000010,
            8'b11111011,
            8'b11111010,
            8'b11111111,
            8'b00000011,
            8'b00000011
        };
    assign keys_wt = '{
            8'b11111110,
            8'b00000000,
            8'b00000010,
            8'b00000010,
            8'b00000010,
            8'b11111111,
            8'b11111000,
            8'b11110110,
            8'b00001010,
            8'b11111111,
            8'b11111010,
            8'b00000001,
            8'b11111111,
            8'b00000010,
            8'b00000001,
            8'b00000100,
            8'b00000111,
            8'b00000110,
            8'b11111011,
            8'b11111110,
            8'b11111101,
            8'b00000101,
            8'b11111100,
            8'b00000011,
            8'b11111011,
            8'b00000001,
            8'b11111111,
            8'b11111110,
            8'b00000011,
            8'b11110101,
            8'b11111010,
            8'b00000001,
            8'b00001000,
            8'b00000101,
            8'b11111110,
            8'b11111111,
            8'b11111110,
            8'b00000111,
            8'b11111111,
            8'b00000101,
            8'b00000100,
            8'b00000010,
            8'b00000001,
            8'b11111110,
            8'b00000000,
            8'b11111100,
            8'b11111110,
            8'b11111111,
            8'b00000010,
            8'b11111101,
            8'b00000010,
            8'b00000010,
            8'b00000000,
            8'b00000100,
            8'b11111110,
            8'b00000011,
            8'b11111110,
            8'b00000000,
            8'b11111110,
            8'b00000001,
            8'b00000110,
            8'b11110110,
            8'b11111000,
            8'b00000000,
            8'b00000000,
            8'b00000011,
            8'b00000110,
            8'b11111110,
            8'b00000111,
            8'b00000100,
            8'b00000001,
            8'b00000011,
            8'b00000001,
            8'b00000001,
            8'b00000101,
            8'b00001001,
            8'b00000011,
            8'b11111100,
            8'b11111000,
            8'b00000000,
            8'b00000100,
            8'b00000101,
            8'b00000001,
            8'b11111100,
            8'b00000100,
            8'b00000011,
            8'b11111111,
            8'b11111110,
            8'b11111111,
            8'b00000000,
            8'b00000001,
            8'b00000001,
            8'b11111101,
            8'b00000000,
            8'b11111000,
            8'b11111110,
            8'b00001101,
            8'b11111111,
            8'b00000101,
            8'b11111011,
            8'b00000100,
            8'b11111101,
            8'b00000000,
            8'b00000001,
            8'b00000000,
            8'b11111111,
            8'b00000010,
            8'b11111111,
            8'b11111110,
            8'b00000000,
            8'b11111010,
            8'b00000011,
            8'b00001001,
            8'b00000011,
            8'b00000100,
            8'b11111111,
            8'b00001100,
            8'b11110111,
            8'b00000000,
            8'b11111010,
            8'b00000001,
            8'b00000111,
            8'b11111100,
            8'b00000000,
            8'b11111100,
            8'b00000110,
            8'b00000110,
            8'b00000011,
            8'b11111110,
            8'b00000001,
            8'b11111110,
            8'b11111110,
            8'b00000000,
            8'b11111111,
            8'b11111111,
            8'b11111110,
            8'b00001000,
            8'b00000101,
            8'b00000000,
            8'b11111111,
            8'b00000100,
            8'b11110010,
            8'b11110100,
            8'b11111110,
            8'b00000111,
            8'b11111101,
            8'b00000001,
            8'b00000000,
            8'b00000010,
            8'b11111110,
            8'b00000100,
            8'b00000001,
            8'b11111110,
            8'b11111110,
            8'b00000100,
            8'b00000101,
            8'b11111101,
            8'b00000100,
            8'b11111000,
            8'b00000001,
            8'b00000101,
            8'b00000011,
            8'b00000001,
            8'b11111101,
            8'b00000000,
            8'b11111101,
            8'b11111101,
            8'b11111101,
            8'b00001000,
            8'b00000101,
            8'b11111100,
            8'b00000010,
            8'b11111110,
            8'b11111111,
            8'b11111101,
            8'b11111110,
            8'b11111100,
            8'b11111001,
            8'b00000011,
            8'b00000011,
            8'b11111101,
            8'b00000011,
            8'b11111110,
            8'b00000011,
            8'b00000011,
            8'b00000011,
            8'b11111111,
            8'b11111100,
            8'b00000111,
            8'b11111001,
            8'b11111000,
            8'b00000011,
            8'b11111110,
            8'b00000001,
            8'b00000001,
            8'b00000010,
            8'b11111100,
            8'b00000100,
            8'b11111111,
            8'b00000011,
            8'b11111000,
            8'b11111111,
            8'b00000011,
            8'b11111011,
            8'b00000000,
            8'b11111000,
            8'b00000001,
            8'b11111001,
            8'b11111111,
            8'b00000001,
            8'b11111011,
            8'b11111111,
            8'b00000010,
            8'b11111010,
            8'b11111100,
            8'b00000000,
            8'b00001001,
            8'b00000011,
            8'b11111100,
            8'b11111100,
            8'b11111011,
            8'b00000001,
            8'b00000010,
            8'b11111110,
            8'b11110111,
            8'b00000010,
            8'b11111100,
            8'b00000010,
            8'b11111111,
            8'b00000010,
            8'b00000000,
            8'b11111011,
            8'b00000001,
            8'b11111101,
            8'b00000100,
            8'b00000000,
            8'b11111011,
            8'b11111111,
            8'b00000011,
            8'b11111100,
            8'b00000001,
            8'b00000100,
            8'b11111110,
            8'b11111100,
            8'b00000110,
            8'b00000010,
            8'b00000000,
            8'b00000001,
            8'b00000001,
            8'b00000001,
            8'b00000001,
            8'b00000001,
            8'b11111101,
            8'b11111011,
            8'b11110111,
            8'b00000010
        };
    assign queries_bs = '{
            8'b11111110,
            8'b11111101,
            8'b00000100,
            8'b00000000,
            8'b00000001,
            8'b00000011,
            8'b00000001,
            8'b00000111,
            8'b00000011,
            8'b00000101,
            8'b00000010,
            8'b11111100,
            8'b11111101,
            8'b00000100,
            8'b11111011,
            8'b00000101
        };
    assign queries_wt = '{
            8'b00000011,
            8'b11111110,
            8'b00000100,
            8'b00000010,
            8'b00000001,
            8'b11111010,
            8'b11111111,
            8'b11111101,
            8'b00000101,
            8'b11111111,
            8'b00000010,
            8'b11111100,
            8'b11111101,
            8'b00000001,
            8'b00000010,
            8'b11111011,
            8'b11111111,
            8'b00000011,
            8'b00000101,
            8'b11111100,
            8'b00000010,
            8'b11111111,
            8'b00000010,
            8'b00000110,
            8'b11111111,
            8'b11111011,
            8'b00000100,
            8'b00001000,
            8'b00000001,
            8'b11111100,
            8'b11110111,
            8'b00000100,
            8'b00000010,
            8'b00000001,
            8'b00000001,
            8'b11111101,
            8'b00000001,
            8'b00000010,
            8'b00000000,
            8'b00000001,
            8'b00000011,
            8'b00000011,
            8'b11111111,
            8'b00000010,
            8'b11111111,
            8'b11111110,
            8'b11111001,
            8'b00000000,
            8'b00000001,
            8'b00000000,
            8'b00000100,
            8'b11111001,
            8'b00000110,
            8'b11111100,
            8'b00000000,
            8'b00000100,
            8'b11111111,
            8'b11111010,
            8'b00000101,
            8'b00001011,
            8'b11111100,
            8'b11111100,
            8'b11111111,
            8'b00000010,
            8'b00000001,
            8'b00000010,
            8'b00000100,
            8'b00000010,
            8'b11111111,
            8'b11111011,
            8'b11111010,
            8'b00000110,
            8'b11111111,
            8'b11111111,
            8'b00000010,
            8'b11111011,
            8'b11111111,
            8'b11111110,
            8'b00000010,
            8'b00001011,
            8'b00000000,
            8'b11111110,
            8'b00000100,
            8'b00000001,
            8'b11111111,
            8'b11111110,
            8'b00000011,
            8'b00000101,
            8'b11111110,
            8'b00000110,
            8'b00000000,
            8'b00000000,
            8'b00000100,
            8'b00000011,
            8'b11111110,
            8'b00000000,
            8'b11111100,
            8'b00000100,
            8'b00000010,
            8'b11111101,
            8'b00000100,
            8'b11111110,
            8'b11111111,
            8'b00000010,
            8'b00000011,
            8'b00000101,
            8'b11111101,
            8'b00000001,
            8'b00000010,
            8'b00000001,
            8'b00000110,
            8'b00000100,
            8'b00000001,
            8'b00000101,
            8'b00000101,
            8'b00000110,
            8'b00000010,
            8'b11111010,
            8'b11111111,
            8'b11111100,
            8'b00000001,
            8'b11111100,
            8'b11110111,
            8'b00000010,
            8'b00000011,
            8'b00000101,
            8'b00001000,
            8'b11111101,
            8'b00000100,
            8'b00000010,
            8'b00000111,
            8'b11111101,
            8'b11111110,
            8'b11111010,
            8'b11111100,
            8'b00000110,
            8'b00000111,
            8'b00000001,
            8'b00001011,
            8'b00000001,
            8'b00000010,
            8'b11111001,
            8'b11111100,
            8'b11111100,
            8'b11111011,
            8'b11111110,
            8'b00000010,
            8'b11111111,
            8'b00000010,
            8'b11111111,
            8'b11111111,
            8'b00000101,
            8'b11111100,
            8'b00000111,
            8'b11111111,
            8'b11111010,
            8'b11111111,
            8'b00000001,
            8'b00000010,
            8'b00000100,
            8'b11111101,
            8'b00000100,
            8'b00000000,
            8'b00000101,
            8'b11111011,
            8'b11111010,
            8'b00000000,
            8'b00000001,
            8'b00000111,
            8'b00000010,
            8'b00000010,
            8'b00000001,
            8'b00000000,
            8'b11111011,
            8'b00000100,
            8'b11111100,
            8'b00000000,
            8'b11111111,
            8'b00000001,
            8'b11111100,
            8'b00000010,
            8'b11111100,
            8'b11111101,
            8'b00000100,
            8'b11111110,
            8'b11111101,
            8'b00000101,
            8'b00000100,
            8'b11111111,
            8'b11111010,
            8'b00000011,
            8'b11111101,
            8'b00000010,
            8'b11111011,
            8'b00000010,
            8'b00000001,
            8'b00000100,
            8'b00000010,
            8'b00000100,
            8'b11111111,
            8'b00000000,
            8'b11111111,
            8'b00000011,
            8'b00000000,
            8'b00000100,
            8'b00000000,
            8'b11111010,
            8'b00000011,
            8'b00000000,
            8'b11111111,
            8'b00000000,
            8'b00001000,
            8'b11111001,
            8'b00000001,
            8'b00000000,
            8'b11111111,
            8'b00001011,
            8'b00000100,
            8'b00000010,
            8'b00000001,
            8'b11111101,
            8'b00000100,
            8'b00000011,
            8'b11110110,
            8'b00000011,
            8'b11111011,
            8'b00000000,
            8'b00000110,
            8'b00000000,
            8'b00001000,
            8'b11111110,
            8'b11111111,
            8'b00000010,
            8'b00000011,
            8'b00000100,
            8'b11111011,
            8'b00000011,
            8'b00000101,
            8'b11111111,
            8'b00000000,
            8'b00000001,
            8'b11111111,
            8'b00000001,
            8'b00000010,
            8'b00000010,
            8'b11111100,
            8'b00000010,
            8'b00000100,
            8'b00000011,
            8'b00000011,
            8'b00000010,
            8'b00000000,
            8'b00000100,
            8'b00000000,
            8'b00000011,
            8'b00000100
        };
    assign values_bs = '{
            8'b11111111,
            8'b11111100,
            8'b00000010,
            8'b11111110,
            8'b00000001,
            8'b11111100,
            8'b11111111,
            8'b00000010,
            8'b11111110,
            8'b11111110,
            8'b00000011,
            8'b00000001,
            8'b11111110,
            8'b00000100,
            8'b00000001,
            8'b11111110
        };
    assign values_wt = '{
            8'b11111110,
            8'b11111110,
            8'b00000010,
            8'b00000101,
            8'b11111110,
            8'b00000110,
            8'b00000001,
            8'b11111101,
            8'b00000001,
            8'b11111010,
            8'b00000110,
            8'b00001101,
            8'b11111100,
            8'b11111100,
            8'b11110111,
            8'b11111001,
            8'b11111000,
            8'b00000001,
            8'b00000101,
            8'b00000111,
            8'b00001011,
            8'b11110010,
            8'b00001001,
            8'b00000001,
            8'b11111010,
            8'b11111111,
            8'b11111111,
            8'b11111101,
            8'b11111111,
            8'b11111010,
            8'b00000101,
            8'b11110001,
            8'b00000001,
            8'b11111100,
            8'b11111011,
            8'b11111010,
            8'b11110101,
            8'b11111101,
            8'b11111010,
            8'b00000011,
            8'b00000010,
            8'b11111000,
            8'b11111001,
            8'b11110100,
            8'b00000111,
            8'b11111011,
            8'b00001000,
            8'b00001101,
            8'b11111010,
            8'b00001000,
            8'b00001000,
            8'b00000101,
            8'b11111111,
            8'b11111100,
            8'b00000110,
            8'b11110111,
            8'b00000000,
            8'b11111010,
            8'b00000110,
            8'b00000100,
            8'b11111100,
            8'b11111110,
            8'b11111011,
            8'b11111010,
            8'b11111010,
            8'b00000101,
            8'b00000101,
            8'b00000000,
            8'b00000010,
            8'b00001000,
            8'b11111111,
            8'b11111111,
            8'b11111101,
            8'b00001100,
            8'b00000010,
            8'b00000100,
            8'b11111010,
            8'b00000001,
            8'b11111101,
            8'b00000100,
            8'b11111100,
            8'b11111001,
            8'b11111011,
            8'b11111010,
            8'b11111110,
            8'b11111011,
            8'b11111111,
            8'b00000011,
            8'b11111110,
            8'b11111010,
            8'b11111001,
            8'b00000000,
            8'b00000100,
            8'b11111101,
            8'b00000110,
            8'b11111011,
            8'b00000010,
            8'b11111100,
            8'b11111000,
            8'b11111001,
            8'b11110111,
            8'b00000111,
            8'b11111011,
            8'b00000011,
            8'b00000101,
            8'b00000100,
            8'b11110111,
            8'b00010000,
            8'b00001001,
            8'b00000010,
            8'b00001000,
            8'b00000110,
            8'b11111011,
            8'b11111110,
            8'b00000001,
            8'b11111101,
            8'b11111111,
            8'b00000000,
            8'b00000011,
            8'b11111101,
            8'b00000000,
            8'b00000110,
            8'b00000010,
            8'b00000010,
            8'b00000000,
            8'b11111101,
            8'b00000110,
            8'b00000001,
            8'b11111100,
            8'b00000011,
            8'b00000001,
            8'b11111111,
            8'b00000100,
            8'b11111101,
            8'b00000011,
            8'b11111100,
            8'b11111110,
            8'b11111100,
            8'b11111101,
            8'b11111001,
            8'b00000000,
            8'b11111100,
            8'b00000000,
            8'b11111111,
            8'b11111000,
            8'b00000001,
            8'b00000010,
            8'b11111101,
            8'b11111001,
            8'b00000001,
            8'b11111110,
            8'b11111011,
            8'b00000110,
            8'b00000001,
            8'b11111100,
            8'b00000010,
            8'b00000000,
            8'b11111100,
            8'b00001101,
            8'b11111111,
            8'b11111011,
            8'b11111101,
            8'b11111000,
            8'b11111100,
            8'b11111111,
            8'b00000011,
            8'b00000010,
            8'b00000101,
            8'b00000100,
            8'b00000101,
            8'b11111100,
            8'b11111000,
            8'b00000100,
            8'b00000111,
            8'b00000101,
            8'b00000010,
            8'b00000111,
            8'b11111100,
            8'b11110111,
            8'b11111111,
            8'b11111001,
            8'b00000010,
            8'b11111001,
            8'b00000111,
            8'b00001001,
            8'b11111010,
            8'b11110110,
            8'b00000000,
            8'b00001000,
            8'b00001000,
            8'b11110111,
            8'b00000110,
            8'b00000011,
            8'b00000110,
            8'b00001011,
            8'b00000010,
            8'b00000110,
            8'b00000110,
            8'b11111111,
            8'b11110101,
            8'b11110111,
            8'b11111110,
            8'b00000111,
            8'b00001000,
            8'b11110111,
            8'b11111100,
            8'b00000001,
            8'b00000100,
            8'b00000100,
            8'b11111101,
            8'b00000011,
            8'b11111111,
            8'b11111011,
            8'b11111110,
            8'b11111110,
            8'b11111101,
            8'b11111110,
            8'b00000001,
            8'b00000011,
            8'b00000000,
            8'b11111101,
            8'b00000001,
            8'b00000010,
            8'b11111110,
            8'b11111101,
            8'b00000001,
            8'b00000000,
            8'b00000010,
            8'b00000101,
            8'b11111101,
            8'b00000100,
            8'b11111100,
            8'b11110100,
            8'b00000001,
            8'b00000101,
            8'b11111110,
            8'b11111111,
            8'b11111101,
            8'b00000110,
            8'b00000000,
            8'b11111100,
            8'b00000100,
            8'b11111111,
            8'b00000101,
            8'b00000000,
            8'b00000001,
            8'b11111111,
            8'b00000010,
            8'b11111111,
            8'b00000100,
            8'b00000100,
            8'b00000001,
            8'b11111100,
            8'b00000000,
            8'b00000111,
            8'b00000001
        };
    assign mlp0_bs = '{
            8'b11111110,
            8'b00000111,
            8'b00000001,
            8'b00000000,
            8'b00000100,
            8'b11111010,
            8'b11111111,
            8'b11111110,
            8'b00000100,
            8'b00000001,
            8'b11111111,
            8'b00000000,
            8'b00000010,
            8'b00000001,
            8'b00000010,
            8'b00000100
        };
    assign mlp0_wt = '{
            8'b00000000,
            8'b11111010,
            8'b11111010,
            8'b00000000,
            8'b00000011,
            8'b00000000,
            8'b00001101,
            8'b00000001,
            8'b11111111,
            8'b00000101,
            8'b11111010,
            8'b11110100,
            8'b00000000,
            8'b00000011,
            8'b00000011,
            8'b00001000,
            8'b11111011,
            8'b00000100,
            8'b00000111,
            8'b00001101,
            8'b00000000,
            8'b11111100,
            8'b11111110,
            8'b11111101,
            8'b11111101,
            8'b11111011,
            8'b11111110,
            8'b00001100,
            8'b00000001,
            8'b00000000,
            8'b00000000,
            8'b00000010,
            8'b00000000,
            8'b11110100,
            8'b00000101,
            8'b00001100,
            8'b00000001,
            8'b11111100,
            8'b00010000,
            8'b00000001,
            8'b00000000,
            8'b11111111,
            8'b11111000,
            8'b00000100,
            8'b11111101,
            8'b00000011,
            8'b00000101,
            8'b00000010,
            8'b00000111,
            8'b11111000,
            8'b00000100,
            8'b00000111,
            8'b00000101,
            8'b00000110,
            8'b11111011,
            8'b00000100,
            8'b11111010,
            8'b00000100,
            8'b00000011,
            8'b11111011,
            8'b00000100,
            8'b11111000,
            8'b11111110,
            8'b00000011,
            8'b11110000,
            8'b00001010,
            8'b11111011,
            8'b00000101,
            8'b00000110,
            8'b11111111,
            8'b11111001,
            8'b11111011,
            8'b11111000,
            8'b11111110,
            8'b00000010,
            8'b00000000,
            8'b00000001,
            8'b11111100,
            8'b11111110,
            8'b00000011,
            8'b00000001,
            8'b11101110,
            8'b00001011,
            8'b00000111,
            8'b00001111,
            8'b11111010,
            8'b00001011,
            8'b00000011,
            8'b00000100,
            8'b00000110,
            8'b11110111,
            8'b11111101,
            8'b11111000,
            8'b00000110,
            8'b00000101,
            8'b11111101,
            8'b00000010,
            8'b11111110,
            8'b11111011,
            8'b11111111,
            8'b00000100,
            8'b00000101,
            8'b00001010,
            8'b00000101,
            8'b00000011,
            8'b00000100,
            8'b11110110,
            8'b00000011,
            8'b11111101,
            8'b00000100,
            8'b00000101,
            8'b00000111,
            8'b00000100,
            8'b00000100,
            8'b00000000,
            8'b00001001,
            8'b00000001,
            8'b00000110,
            8'b00001100,
            8'b11111111,
            8'b00000110,
            8'b00000101,
            8'b11111011,
            8'b11110001,
            8'b11111100,
            8'b00000101,
            8'b00000111,
            8'b11110100,
            8'b11111110,
            8'b00000010,
            8'b00000000,
            8'b00000100,
            8'b11111100,
            8'b11111100,
            8'b11111000,
            8'b00000001,
            8'b11111110,
            8'b00000100,
            8'b11111001,
            8'b00001100,
            8'b11111111,
            8'b11111110,
            8'b00000011,
            8'b00000001,
            8'b00000100,
            8'b11111011,
            8'b00000000,
            8'b00000110,
            8'b00000110,
            8'b11111011,
            8'b00000001,
            8'b00000011,
            8'b00000001,
            8'b00000100,
            8'b00000001,
            8'b00001010,
            8'b11111100,
            8'b00000001,
            8'b00000011,
            8'b00000001,
            8'b11111111,
            8'b11110101,
            8'b11110110,
            8'b11111010,
            8'b11110100,
            8'b11111110,
            8'b00000111,
            8'b00000101,
            8'b00000001,
            8'b11111011,
            8'b11111010,
            8'b00000001,
            8'b11111100,
            8'b00000011,
            8'b00000011,
            8'b11111110,
            8'b00000001,
            8'b11111101,
            8'b11111001,
            8'b11111101,
            8'b11110111,
            8'b11111110,
            8'b00000011,
            8'b00000001,
            8'b00000011,
            8'b11111101,
            8'b11111010,
            8'b00000101,
            8'b11111101,
            8'b00000010,
            8'b00000101,
            8'b00001001,
            8'b11111101,
            8'b00000111,
            8'b11111001,
            8'b00001010,
            8'b00000100,
            8'b00001010,
            8'b00000100,
            8'b11110000,
            8'b11111110,
            8'b00000001,
            8'b00000110,
            8'b00001000,
            8'b00000001,
            8'b11111111,
            8'b11111110,
            8'b00000000,
            8'b00000110,
            8'b00000001,
            8'b11111001,
            8'b11111110,
            8'b00001000,
            8'b00000000,
            8'b00000000,
            8'b00000000,
            8'b00000011,
            8'b00001001,
            8'b11110111,
            8'b00001001,
            8'b11111100,
            8'b11111111,
            8'b00000101,
            8'b00000111,
            8'b11111100,
            8'b00000011,
            8'b11111010,
            8'b11111111,
            8'b00000000,
            8'b00000111,
            8'b11110011,
            8'b00000011,
            8'b11111010,
            8'b11110000,
            8'b00000001,
            8'b00001011,
            8'b00000000,
            8'b11111011,
            8'b11111011,
            8'b00000001,
            8'b11110111,
            8'b11111011,
            8'b00000001,
            8'b11110010,
            8'b00000110,
            8'b00001100,
            8'b11111111,
            8'b00000101,
            8'b00000001,
            8'b00000100,
            8'b11111110,
            8'b11111010,
            8'b11111110,
            8'b11111110,
            8'b00000001,
            8'b00000100
        };
    assign mlp1_bs = '{
            8'b11111110,
            8'b11111111,
            8'b00000001,
            8'b11111111,
            8'b11111010,
            8'b00000001,
            8'b00000011,
            8'b00000010,
            8'b00000000,
            8'b11111111,
            8'b00000000,
            8'b11111111,
            8'b00000000,
            8'b11111111,
            8'b11111101,
            8'b11111111
        };
    assign mlp1_wt = '{
            8'b00000001,
            8'b11111110,
            8'b00000011,
            8'b00000001,
            8'b11110111,
            8'b00000100,
            8'b00000010,
            8'b11111010,
            8'b00000010,
            8'b00001010,
            8'b11111100,
            8'b11111010,
            8'b00000111,
            8'b11111111,
            8'b00000010,
            8'b00000011,
            8'b11111111,
            8'b11111101,
            8'b11110111,
            8'b11111010,
            8'b00001101,
            8'b00000101,
            8'b00000011,
            8'b11111100,
            8'b11111111,
            8'b11111001,
            8'b00000011,
            8'b00000010,
            8'b00000001,
            8'b00000101,
            8'b11111111,
            8'b11111010,
            8'b00000111,
            8'b11111110,
            8'b11111100,
            8'b00000100,
            8'b11111001,
            8'b00000011,
            8'b00000010,
            8'b11111100,
            8'b11111110,
            8'b11111011,
            8'b11111011,
            8'b00000100,
            8'b11110110,
            8'b00000011,
            8'b00000101,
            8'b11111000,
            8'b11111011,
            8'b00000111,
            8'b00000011,
            8'b11111011,
            8'b00000001,
            8'b00000001,
            8'b11111101,
            8'b00001000,
            8'b00000000,
            8'b00000001,
            8'b11111101,
            8'b11111110,
            8'b00000001,
            8'b11111100,
            8'b00000101,
            8'b00000001,
            8'b00000111,
            8'b11110111,
            8'b00000000,
            8'b00000111,
            8'b11110110,
            8'b00000001,
            8'b00000011,
            8'b11111001,
            8'b11111111,
            8'b00000010,
            8'b11111100,
            8'b00000001,
            8'b11111010,
            8'b00000100,
            8'b00000011,
            8'b11111110,
            8'b00000001,
            8'b00000011,
            8'b11111100,
            8'b11111100,
            8'b00000010,
            8'b00000110,
            8'b11111110,
            8'b00000010,
            8'b11111110,
            8'b11111001,
            8'b11111100,
            8'b11111111,
            8'b11111101,
            8'b00000010,
            8'b00000101,
            8'b11111011,
            8'b11111110,
            8'b00000010,
            8'b00000011,
            8'b11111111,
            8'b00000011,
            8'b11111001,
            8'b00000000,
            8'b00000010,
            8'b00000101,
            8'b00000010,
            8'b00000110,
            8'b11111110,
            8'b00000001,
            8'b11111100,
            8'b11111010,
            8'b00000111,
            8'b00000110,
            8'b11111010,
            8'b00000001,
            8'b00001010,
            8'b11111101,
            8'b11111001,
            8'b00000111,
            8'b11110110,
            8'b11111100,
            8'b00000001,
            8'b00000101,
            8'b00000011,
            8'b11111001,
            8'b00000101,
            8'b11111010,
            8'b11111101,
            8'b00000100,
            8'b11111110,
            8'b00000010,
            8'b00000100,
            8'b11111111,
            8'b11110110,
            8'b00000110,
            8'b11111010,
            8'b11111110,
            8'b11111110,
            8'b00001001,
            8'b00000010,
            8'b11111001,
            8'b00000100,
            8'b11111010,
            8'b00000001,
            8'b00000101,
            8'b11111001,
            8'b00000000,
            8'b00000100,
            8'b00000010,
            8'b11111011,
            8'b00000001,
            8'b11111000,
            8'b00000010,
            8'b00000001,
            8'b00000101,
            8'b00000111,
            8'b11111111,
            8'b00000011,
            8'b11111001,
            8'b00000010,
            8'b11111100,
            8'b00000110,
            8'b00000000,
            8'b11111111,
            8'b11111111,
            8'b00000011,
            8'b11111111,
            8'b00000111,
            8'b11111110,
            8'b11111111,
            8'b11111011,
            8'b11111110,
            8'b11111101,
            8'b11111110,
            8'b00000111,
            8'b11111100,
            8'b11111111,
            8'b11111101,
            8'b11111111,
            8'b11111111,
            8'b11111010,
            8'b00000100,
            8'b00000010,
            8'b11111100,
            8'b00000011,
            8'b00000110,
            8'b11111110,
            8'b11111111,
            8'b00001101,
            8'b11111100,
            8'b00000001,
            8'b00000001,
            8'b11111111,
            8'b00000101,
            8'b11111101,
            8'b11111001,
            8'b00000010,
            8'b00001010,
            8'b11111001,
            8'b00000111,
            8'b00000100,
            8'b11111101,
            8'b11111011,
            8'b11111010,
            8'b00000111,
            8'b11111110,
            8'b00000100,
            8'b00000011,
            8'b00000011,
            8'b11111010,
            8'b00000100,
            8'b00001001,
            8'b11111100,
            8'b11111000,
            8'b00000010,
            8'b11111011,
            8'b00000001,
            8'b11111111,
            8'b00000101,
            8'b00000101,
            8'b11111010,
            8'b00000010,
            8'b11111000,
            8'b00000100,
            8'b00000011,
            8'b11110111,
            8'b11111011,
            8'b00000010,
            8'b11111011,
            8'b00000010,
            8'b00000110,
            8'b11110110,
            8'b00000000,
            8'b11111111,
            8'b11111111,
            8'b00000110,
            8'b00000101,
            8'b00000011,
            8'b11111101,
            8'b11111101,
            8'b00000000,
            8'b00000100,
            8'b00001000,
            8'b00000111,
            8'b11111011,
            8'b11111111,
            8'b00000011,
            8'b00000011,
            8'b00000001,
            8'b11111101,
            8'b11111010,
            8'b11111101,
            8'b11110001,
            8'b11111011,
            8'b00000011,
            8'b00000001
        };
    assign ps_wt = '{
            8'b00001100,
            8'b00000000,
            8'b11101000,
            8'b11101110,
            8'b00000111,
            8'b11111001,
            8'b00001100,
            8'b00011100,
            8'b00011001,
            8'b11111111,
            8'b00001010,
            8'b00001010,
            8'b11100111,
            8'b00001000,
            8'b11101001,
            8'b11110001,
            8'b00010001,
            8'b11110111,
            8'b11111100,
            8'b00001100,
            8'b00000110,
            8'b11011011,
            8'b11111011,
            8'b11111011,
            8'b11110000,
            8'b11100100,
            8'b11111000,
            8'b00001000,
            8'b00001001,
            8'b00000100,
            8'b11110101,
            8'b00000001,
            8'b00000011,
            8'b11100001,
            8'b00101010,
            8'b11111001,
            8'b11101000,
            8'b11110000,
            8'b11011100,
            8'b00000101,
            8'b11111001,
            8'b11100101,
            8'b11110110,
            8'b11110011,
            8'b00001101,
            8'b00010111,
            8'b00100000,
            8'b11101010,
            8'b00001100,
            8'b00011101,
            8'b00010110,
            8'b00000100,
            8'b11111011,
            8'b00000101,
            8'b11101010,
            8'b00010000,
            8'b00000100,
            8'b00001100,
            8'b00100011,
            8'b00010000,
            8'b11110000,
            8'b00000000,
            8'b00000110,
            8'b00010110,
            8'b00001000,
            8'b11110010,
            8'b00000011,
            8'b00000100,
            8'b11100100,
            8'b00010010,
            8'b00001100,
            8'b00000001,
            8'b00000001,
            8'b00000001,
            8'b00001100,
            8'b00001101,
            8'b00010100,
            8'b00001010,
            8'b11100010,
            8'b11110111,
            8'b11100011,
            8'b00000000,
            8'b11111100,
            8'b11111111,
            8'b00010111,
            8'b11011000,
            8'b00100010,
            8'b00110100,
            8'b11111000,
            8'b00000101,
            8'b00000110,
            8'b11101011,
            8'b00001001,
            8'b00001001,
            8'b00010000,
            8'b11111110,
            8'b00000010,
            8'b00010100,
            8'b00011001,
            8'b00001110,
            8'b00010000,
            8'b11110111,
            8'b11010111,
            8'b00000101,
            8'b00010101,
            8'b00100001,
            8'b11101101,
            8'b00001101,
            8'b00001111,
            8'b11110110,
            8'b00000000,
            8'b00010111,
            8'b11110001,
            8'b11101110,
            8'b11110101,
            8'b00010110,
            8'b00000100,
            8'b11111001,
            8'b00000000,
            8'b11111101,
            8'b00011010,
            8'b00010100,
            8'b11111111,
            8'b00000000,
            8'b00000001,
            8'b00010000,
            8'b00011001,
            8'b11111000,
            8'b00010100,
            8'b11111010,
            8'b00001000,
            8'b11110010,
            8'b00001000,
            8'b11101111,
            8'b11111011,
            8'b11110001,
            8'b00110001,
            8'b00010101,
            8'b00001011,
            8'b00000001,
            8'b11111101,
            8'b00011000,
            8'b11011111,
            8'b00100000,
            8'b11111111,
            8'b11111101,
            8'b00000001,
            8'b00010100,
            8'b11111011,
            8'b11101100,
            8'b11011010,
            8'b11110100,
            8'b00000010,
            8'b00010011,
            8'b11100101,
            8'b11100011,
            8'b00000011,
            8'b11111100,
            8'b11111001,
            8'b00001000,
            8'b11011101,
            8'b11100100,
            8'b11110011,
            8'b11101111,
            8'b11111100,
            8'b11110001,
            8'b11110000,
            8'b00011000,
            8'b11110110,
            8'b11100110,
            8'b11100100,
            8'b00000011,
            8'b00011100,
            8'b11101111,
            8'b00000010,
            8'b00010101,
            8'b11111010,
            8'b00010001,
            8'b11110011,
            8'b11111111,
            8'b11011100,
            8'b00011011,
            8'b11111101,
            8'b00010011,
            8'b11111111,
            8'b00001101,
            8'b11110001,
            8'b11101110,
            8'b11111110,
            8'b00010100,
            8'b00000011,
            8'b11110101,
            8'b11110110,
            8'b00010111,
            8'b11101101,
            8'b11110111,
            8'b00000110,
            8'b00011000,
            8'b00010011,
            8'b11110000,
            8'b11110010,
            8'b11111010,
            8'b11101001,
            8'b00000111,
            8'b11101100,
            8'b00000001,
            8'b11111111,
            8'b00010001,
            8'b11110101,
            8'b11111101,
            8'b00100000,
            8'b11100010,
            8'b00001010,
            8'b11101111,
            8'b00010000,
            8'b11111111,
            8'b11101001,
            8'b00011001,
            8'b11101001,
            8'b00001100,
            8'b11110011,
            8'b00001001,
            8'b11110011,
            8'b00010011,
            8'b11110010,
            8'b11110001,
            8'b11110100,
            8'b00010010,
            8'b11100101,
            8'b00000100,
            8'b00010101,
            8'b11110010,
            8'b11111110,
            8'b00010011,
            8'b11110110,
            8'b11100111,
            8'b00001111,
            8'b00011111,
            8'b11101100,
            8'b11100111,
            8'b00100001,
            8'b00101111,
            8'b11011110,
            8'b00011001,
            8'b11111000,
            8'b00000011,
            8'b00010110,
            8'b00001000,
            8'b00001111,
            8'b00011000,
            8'b11111000,
            8'b11110100,
            8'b00011001,
            8'b11111011,
            8'b00011010,
            8'b00001011
        };



    // Output logic
    always_comb begin
        case (addr)
            8'h01:   data_o = classifier_bs;
            8'h02:   data_o = classifier_wt;
            8'h03:   data_o = embedding_bs;
            8'h04:   data_o = embedding_wt;
            8'h05:   data_o = cls_token_wt;
            8'h06:   data_o = final_bs;
            8'h07:   data_o = final_wt;
            8'h08:   data_o = keys_bs;
            8'h09:   data_o = keys_wt;
            8'h0A:   data_o = queries_bs;
            8'h0B:   data_o = queries_wt;
            8'h0C:   data_o = values_bs;
            8'h0D:   data_o = values_wt;
            8'h0E:   data_o = mlp0_bs;
            8'h0F:   data_o = mlp0_wt;
            8'h10:   data_o = mlp1_bs;
            8'h11:   data_o = mlp1_wt;
            8'h12:   data_o = ps_wt;
            default: data_o = '{default: '0};
        endcase
    end

endmodule
