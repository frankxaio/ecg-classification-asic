module lut_module #(
    parameter ADDR_WIDTH = 8,
    parameter DATA_WIDTH = 8
) (
    input                         clk,
    input                         rst,
    input                         start,
    input        [ADDR_WIDTH-1:0] addr,
    output logic [DATA_WIDTH-1:0] data_o,
    output logic                  done
);

    localparam CLASSIFIER_BS_CNT = 6;
    localparam CLASSIFIER_WT_CNT = 96;
    localparam EMBEDDING_BS_CNT = 16;
    localparam EMBEDDING_WT_CNT = 16;
    localparam CLS_TOKEN_WT_CNT = 16;
    localparam FINAL_BS_CNT = 16;
    localparam FINAL_WT_CNT = 256;
    localparam KEYS_BS_CNT = 16;
    localparam KEYS_WT_CNT = 256;
    localparam QUERIES_BS_CNT = 16;
    localparam QUERIES_WT_CNT = 256;
    localparam VALUES_BS_CNT = 16;
    localparam VALUES_WT_CNT = 256;
    localparam MLP0_BS_CNT = 16;
    localparam MLP0_WT_CNT = 256;
    localparam MLP1_BS_CNT = 16;
    localparam MLP1_WT_CNT = 256;
    localparam PS_WT_CNT = 256;

    // Define the memory arrays for each file
    logic [DATA_WIDTH-1:0] classifier_bs[0:5];
    logic [DATA_WIDTH-1:0] classifier_wt[0:95];
    logic [DATA_WIDTH-1:0] embedding_bs[0:15];
    logic [DATA_WIDTH-1:0] embedding_wt[0:15];
    logic [DATA_WIDTH-1:0] cls_token_wt[0:15];
    logic [DATA_WIDTH-1:0] final_bs[0:15];
    logic [DATA_WIDTH-1:0] final_wt[0:255];
    logic [DATA_WIDTH-1:0] keys_bs[0:15];
    logic [DATA_WIDTH-1:0] keys_wt[0:255];
    logic [DATA_WIDTH-1:0] queries_bs[0:15];
    logic [DATA_WIDTH-1:0] queries_wt[0:255];
    logic [DATA_WIDTH-1:0] values_bs[0:15];
    logic [DATA_WIDTH-1:0] values_wt[0:255];
    logic [DATA_WIDTH-1:0] mlp0_bs[0:15];
    logic [DATA_WIDTH-1:0] mlp0_wt[0:255];
    logic [DATA_WIDTH-1:0] mlp1_bs[0:15];
    logic [DATA_WIDTH-1:0] mlp1_wt[0:255];
    logic [DATA_WIDTH-1:0] ps_wt[0:255];

    // Array index register
    logic [$clog2(256):0] array_index, array_index_ns;
    logic [DATA_WIDTH-1:0] data;


    //LUT DATA
    assign classifier_bs = {
        8'b00000100, 8'b11111111, 8'b00000000, 8'b11111001, 8'b00000000, 8'b11111010
    };
    assign classifier_wt = {
        8'b00000100,
        8'b11111011,
        8'b11111001,
        8'b11111010,
        8'b00000011,
        8'b11111000,
        8'b00001000,
        8'b00000111,
        8'b00000110,
        8'b00001000,
        8'b11111010,
        8'b00000000,
        8'b11111001,
        8'b00001000,
        8'b00000001,
        8'b00000000,
        8'b00001001,
        8'b00010010,
        8'b00001110,
        8'b11110101,
        8'b00001100,
        8'b00000100,
        8'b11101100,
        8'b00000010,
        8'b00000000,
        8'b00000011,
        8'b11110111,
        8'b00010110,
        8'b11111100,
        8'b11111111,
        8'b00001111,
        8'b11101101,
        8'b00001010,
        8'b11101101,
        8'b11111111,
        8'b00001110,
        8'b00000001,
        8'b00000001,
        8'b11111011,
        8'b11111011,
        8'b11110101,
        8'b11111010,
        8'b00001010,
        8'b00001110,
        8'b00000111,
        8'b11111000,
        8'b11111001,
        8'b00001011,
        8'b11111111,
        8'b11011000,
        8'b00001101,
        8'b00001101,
        8'b00001110,
        8'b00000100,
        8'b00000010,
        8'b11111110,
        8'b11111110,
        8'b11111010,
        8'b00000001,
        8'b11111101,
        8'b11111001,
        8'b00000010,
        8'b00000100,
        8'b00000010,
        8'b11110110,
        8'b00010010,
        8'b11101111,
        8'b00010100,
        8'b11101111,
        8'b00001111,
        8'b00000111,
        8'b11110011,
        8'b11110110,
        8'b11111001,
        8'b00001101,
        8'b11110001,
        8'b00001100,
        8'b11110001,
        8'b11110010,
        8'b11111010,
        8'b11111100,
        8'b00000111,
        8'b00001111,
        8'b11110110,
        8'b00000101,
        8'b00000110,
        8'b11111011,
        8'b00000110,
        8'b00000110,
        8'b00000011,
        8'b00000010,
        8'b11101101,
        8'b11111001,
        8'b00000011,
        8'b00000000,
        8'b00000101
    };
    assign embedding_bs = {
        8'b11111010,
        8'b00010000,
        8'b11110010,
        8'b00001011,
        8'b11111101,
        8'b00000010,
        8'b11110101,
        8'b00001111,
        8'b00010001,
        8'b11111010,
        8'b00000000,
        8'b11110001,
        8'b00000111,
        8'b00001010,
        8'b00010001,
        8'b00000100
    };
    assign embedding_wt = {
        8'b00001100,
        8'b11110001,
        8'b00001101,
        8'b11100100,
        8'b00000001,
        8'b00000101,
        8'b00000100,
        8'b00010110,
        8'b11101110,
        8'b11111101,
        8'b11111010,
        8'b11111101,
        8'b00010011,
        8'b11101000,
        8'b11011111,
        8'b00011011
    };
    assign cls_token_wt = {
        8'b00000111,
        8'b00001111,
        8'b00000101,
        8'b11101001,
        8'b00001101,
        8'b00000100,
        8'b11111110,
        8'b00000011,
        8'b11111111,
        8'b11101101,
        8'b00010100,
        8'b00000011,
        8'b00000001,
        8'b00000110,
        8'b00001100,
        8'b00000110
    };
    assign final_bs = {
        8'b00000011,
        8'b00000011,
        8'b11111100,
        8'b11111110,
        8'b11111101,
        8'b00000000,
        8'b11111110,
        8'b00000010,
        8'b00000110,
        8'b00000100,
        8'b00000010,
        8'b00000010,
        8'b11111111,
        8'b00000101,
        8'b00000010,
        8'b00000000
    };
    assign final_wt = {
        8'b11111110,
        8'b00000010,
        8'b00000011,
        8'b00000110,
        8'b00000100,
        8'b00000111,
        8'b11111111,
        8'b11111111,
        8'b00000000,
        8'b00000100,
        8'b00000110,
        8'b11111111,
        8'b11111100,
        8'b00000100,
        8'b11111011,
        8'b00000101,
        8'b00000100,
        8'b00000000,
        8'b11111111,
        8'b00000111,
        8'b00000000,
        8'b11111101,
        8'b11111001,
        8'b00000101,
        8'b11111111,
        8'b11111011,
        8'b11111110,
        8'b00001000,
        8'b00000001,
        8'b00000011,
        8'b11111100,
        8'b00000000,
        8'b11111101,
        8'b11111110,
        8'b00000000,
        8'b00000011,
        8'b11111101,
        8'b00000010,
        8'b00000001,
        8'b11111101,
        8'b11111111,
        8'b00001110,
        8'b00000000,
        8'b11111101,
        8'b11111110,
        8'b00000100,
        8'b00000010,
        8'b00000001,
        8'b11111011,
        8'b11111110,
        8'b11111101,
        8'b11111101,
        8'b00000011,
        8'b00000000,
        8'b11111111,
        8'b00000000,
        8'b11111110,
        8'b00000011,
        8'b11111111,
        8'b11111111,
        8'b00000001,
        8'b00000010,
        8'b00000100,
        8'b00000101,
        8'b00000011,
        8'b00000011,
        8'b00000010,
        8'b11110111,
        8'b11111001,
        8'b00000010,
        8'b11111100,
        8'b11111011,
        8'b11111111,
        8'b00000111,
        8'b00000011,
        8'b11111100,
        8'b00000010,
        8'b11111100,
        8'b00000101,
        8'b00001110,
        8'b00000101,
        8'b00000000,
        8'b00000001,
        8'b11111100,
        8'b11101111,
        8'b00010111,
        8'b11101111,
        8'b11111101,
        8'b00000101,
        8'b00000100,
        8'b00000010,
        8'b00010001,
        8'b11111101,
        8'b00000100,
        8'b11111111,
        8'b00001010,
        8'b11111001,
        8'b00000011,
        8'b00000000,
        8'b00000011,
        8'b00000110,
        8'b00000001,
        8'b00000000,
        8'b11111100,
        8'b11111100,
        8'b00000001,
        8'b00000001,
        8'b00001001,
        8'b00000001,
        8'b11111011,
        8'b00000111,
        8'b11111011,
        8'b11111100,
        8'b00000100,
        8'b00000101,
        8'b00000101,
        8'b00000000,
        8'b00000001,
        8'b00000001,
        8'b11111110,
        8'b00000011,
        8'b00000000,
        8'b00000010,
        8'b00000010,
        8'b00000001,
        8'b00000001,
        8'b11111101,
        8'b11111011,
        8'b00000001,
        8'b00000101,
        8'b00001101,
        8'b00000100,
        8'b00000111,
        8'b00000101,
        8'b00001001,
        8'b11110110,
        8'b11111100,
        8'b00000111,
        8'b00001111,
        8'b00010100,
        8'b11110100,
        8'b11111011,
        8'b11111010,
        8'b11111001,
        8'b00000001,
        8'b00000111,
        8'b00000110,
        8'b00000001,
        8'b00000111,
        8'b00000101,
        8'b11111110,
        8'b00000000,
        8'b11111010,
        8'b00000110,
        8'b00000100,
        8'b00000000,
        8'b11111011,
        8'b00000001,
        8'b00000011,
        8'b00001000,
        8'b00000011,
        8'b11111100,
        8'b11111011,
        8'b11111000,
        8'b00000001,
        8'b00000111,
        8'b00000101,
        8'b00000101,
        8'b00000000,
        8'b00001001,
        8'b00000001,
        8'b11111100,
        8'b00000101,
        8'b00000011,
        8'b11111110,
        8'b00000000,
        8'b00000100,
        8'b00000010,
        8'b11111100,
        8'b11111101,
        8'b00000101,
        8'b11111011,
        8'b00000000,
        8'b00000001,
        8'b11111011,
        8'b11111011,
        8'b11111100,
        8'b11110001,
        8'b00000101,
        8'b11111101,
        8'b00000000,
        8'b00000101,
        8'b11111111,
        8'b11110111,
        8'b11101110,
        8'b11110111,
        8'b11111111,
        8'b00000101,
        8'b11110110,
        8'b00010101,
        8'b00001011,
        8'b00001010,
        8'b11110010,
        8'b11111001,
        8'b00001101,
        8'b00001100,
        8'b00000010,
        8'b00000111,
        8'b11111111,
        8'b00000101,
        8'b00001110,
        8'b00000100,
        8'b00000101,
        8'b11111101,
        8'b00001001,
        8'b11110110,
        8'b11110010,
        8'b00000001,
        8'b00001100,
        8'b00001000,
        8'b11110011,
        8'b11111000,
        8'b11111111,
        8'b11110100,
        8'b11111111,
        8'b00000101,
        8'b00001111,
        8'b00000110,
        8'b11111111,
        8'b11111110,
        8'b00000101,
        8'b11110100,
        8'b11111010,
        8'b11111111,
        8'b00001000,
        8'b00000100,
        8'b11111001,
        8'b11111001,
        8'b11111110,
        8'b00000001,
        8'b11111110,
        8'b00000001,
        8'b00000011,
        8'b00000011,
        8'b11111101,
        8'b11111111,
        8'b11111100,
        8'b11111110,
        8'b00000001,
        8'b11111000,
        8'b11111101,
        8'b00000000,
        8'b00000010,
        8'b11111110,
        8'b00000010,
        8'b00000101
    };
    assign keys_bs = {
        8'b00000100,
        8'b11110111,
        8'b11111111,
        8'b11110011,
        8'b00000001,
        8'b11111111,
        8'b00000001,
        8'b00000001,
        8'b11111100,
        8'b00001001,
        8'b00000010,
        8'b11111011,
        8'b11111010,
        8'b11111111,
        8'b00000011,
        8'b00000011
    };
    assign keys_wt = {
        8'b11111110,
        8'b00000000,
        8'b00000010,
        8'b00000010,
        8'b00000010,
        8'b11111111,
        8'b11111000,
        8'b11110110,
        8'b00001010,
        8'b11111111,
        8'b11111010,
        8'b00000001,
        8'b11111111,
        8'b00000010,
        8'b00000001,
        8'b00000100,
        8'b00000111,
        8'b00000110,
        8'b11111011,
        8'b11111110,
        8'b11111101,
        8'b00000101,
        8'b11111100,
        8'b00000011,
        8'b11111011,
        8'b00000001,
        8'b11111111,
        8'b11111110,
        8'b00000011,
        8'b11110101,
        8'b11111010,
        8'b00000001,
        8'b00001000,
        8'b00000101,
        8'b11111110,
        8'b11111111,
        8'b11111110,
        8'b00000111,
        8'b11111111,
        8'b00000101,
        8'b00000100,
        8'b00000010,
        8'b00000001,
        8'b11111110,
        8'b00000000,
        8'b11111100,
        8'b11111110,
        8'b11111111,
        8'b00000010,
        8'b11111101,
        8'b00000010,
        8'b00000010,
        8'b00000000,
        8'b00000100,
        8'b11111110,
        8'b00000011,
        8'b11111110,
        8'b00000000,
        8'b11111110,
        8'b00000001,
        8'b00000110,
        8'b11110110,
        8'b11111000,
        8'b00000000,
        8'b00000000,
        8'b00000011,
        8'b00000110,
        8'b11111110,
        8'b00000111,
        8'b00000100,
        8'b00000001,
        8'b00000011,
        8'b00000001,
        8'b00000001,
        8'b00000101,
        8'b00001001,
        8'b00000011,
        8'b11111100,
        8'b11111000,
        8'b00000000,
        8'b00000100,
        8'b00000101,
        8'b00000001,
        8'b11111100,
        8'b00000100,
        8'b00000011,
        8'b11111111,
        8'b11111110,
        8'b11111111,
        8'b00000000,
        8'b00000001,
        8'b00000001,
        8'b11111101,
        8'b00000000,
        8'b11111000,
        8'b11111110,
        8'b00001101,
        8'b11111111,
        8'b00000101,
        8'b11111011,
        8'b00000100,
        8'b11111101,
        8'b00000000,
        8'b00000001,
        8'b00000000,
        8'b11111111,
        8'b00000010,
        8'b11111111,
        8'b11111110,
        8'b00000000,
        8'b11111010,
        8'b00000011,
        8'b00001001,
        8'b00000011,
        8'b00000100,
        8'b11111111,
        8'b00001100,
        8'b11110111,
        8'b00000000,
        8'b11111010,
        8'b00000001,
        8'b00000111,
        8'b11111100,
        8'b00000000,
        8'b11111100,
        8'b00000110,
        8'b00000110,
        8'b00000011,
        8'b11111110,
        8'b00000001,
        8'b11111110,
        8'b11111110,
        8'b00000000,
        8'b11111111,
        8'b11111111,
        8'b11111110,
        8'b00001000,
        8'b00000101,
        8'b00000000,
        8'b11111111,
        8'b00000100,
        8'b11110010,
        8'b11110100,
        8'b11111110,
        8'b00000111,
        8'b11111101,
        8'b00000001,
        8'b00000000,
        8'b00000010,
        8'b11111110,
        8'b00000100,
        8'b00000001,
        8'b11111110,
        8'b11111110,
        8'b00000100,
        8'b00000101,
        8'b11111101,
        8'b00000100,
        8'b11111000,
        8'b00000001,
        8'b00000101,
        8'b00000011,
        8'b00000001,
        8'b11111101,
        8'b00000000,
        8'b11111101,
        8'b11111101,
        8'b11111101,
        8'b00001000,
        8'b00000101,
        8'b11111100,
        8'b00000010,
        8'b11111110,
        8'b11111111,
        8'b11111101,
        8'b11111110,
        8'b11111100,
        8'b11111001,
        8'b00000011,
        8'b00000011,
        8'b11111101,
        8'b00000011,
        8'b11111110,
        8'b00000011,
        8'b00000011,
        8'b00000011,
        8'b11111111,
        8'b11111100,
        8'b00000111,
        8'b11111001,
        8'b11111000,
        8'b00000011,
        8'b11111110,
        8'b00000001,
        8'b00000001,
        8'b00000010,
        8'b11111100,
        8'b00000100,
        8'b11111111,
        8'b00000011,
        8'b11111000,
        8'b11111111,
        8'b00000011,
        8'b11111011,
        8'b00000000,
        8'b11111000,
        8'b00000001,
        8'b11111001,
        8'b11111111,
        8'b00000001,
        8'b11111011,
        8'b11111111,
        8'b00000010,
        8'b11111010,
        8'b11111100,
        8'b00000000,
        8'b00001001,
        8'b00000011,
        8'b11111100,
        8'b11111100,
        8'b11111011,
        8'b00000001,
        8'b00000010,
        8'b11111110,
        8'b11110111,
        8'b00000010,
        8'b11111100,
        8'b00000010,
        8'b11111111,
        8'b00000010,
        8'b00000000,
        8'b11111011,
        8'b00000001,
        8'b11111101,
        8'b00000100,
        8'b00000000,
        8'b11111011,
        8'b11111111,
        8'b00000011,
        8'b11111100,
        8'b00000001,
        8'b00000100,
        8'b11111110,
        8'b11111100,
        8'b00000110,
        8'b00000010,
        8'b00000000,
        8'b00000001,
        8'b00000001,
        8'b00000001,
        8'b00000001,
        8'b00000001,
        8'b11111101,
        8'b11111011,
        8'b11110111,
        8'b00000010
    };
    assign queries_bs = {
        8'b11111110,
        8'b11111101,
        8'b00000100,
        8'b00000000,
        8'b00000001,
        8'b00000011,
        8'b00000001,
        8'b00000111,
        8'b00000011,
        8'b00000101,
        8'b00000010,
        8'b11111100,
        8'b11111101,
        8'b00000100,
        8'b11111011,
        8'b00000101
    };
    assign queries_wt = {
        8'b00000011,
        8'b11111110,
        8'b00000100,
        8'b00000010,
        8'b00000001,
        8'b11111010,
        8'b11111111,
        8'b11111101,
        8'b00000101,
        8'b11111111,
        8'b00000010,
        8'b11111100,
        8'b11111101,
        8'b00000001,
        8'b00000010,
        8'b11111011,
        8'b11111111,
        8'b00000011,
        8'b00000101,
        8'b11111100,
        8'b00000010,
        8'b11111111,
        8'b00000010,
        8'b00000110,
        8'b11111111,
        8'b11111011,
        8'b00000100,
        8'b00001000,
        8'b00000001,
        8'b11111100,
        8'b11110111,
        8'b00000100,
        8'b00000010,
        8'b00000001,
        8'b00000001,
        8'b11111101,
        8'b00000001,
        8'b00000010,
        8'b00000000,
        8'b00000001,
        8'b00000011,
        8'b00000011,
        8'b11111111,
        8'b00000010,
        8'b11111111,
        8'b11111110,
        8'b11111001,
        8'b00000000,
        8'b00000001,
        8'b00000000,
        8'b00000100,
        8'b11111001,
        8'b00000110,
        8'b11111100,
        8'b00000000,
        8'b00000100,
        8'b11111111,
        8'b11111010,
        8'b00000101,
        8'b00001011,
        8'b11111100,
        8'b11111100,
        8'b11111111,
        8'b00000010,
        8'b00000001,
        8'b00000010,
        8'b00000100,
        8'b00000010,
        8'b11111111,
        8'b11111011,
        8'b11111010,
        8'b00000110,
        8'b11111111,
        8'b11111111,
        8'b00000010,
        8'b11111011,
        8'b11111111,
        8'b11111110,
        8'b00000010,
        8'b00001011,
        8'b00000000,
        8'b11111110,
        8'b00000100,
        8'b00000001,
        8'b11111111,
        8'b11111110,
        8'b00000011,
        8'b00000101,
        8'b11111110,
        8'b00000110,
        8'b00000000,
        8'b00000000,
        8'b00000100,
        8'b00000011,
        8'b11111110,
        8'b00000000,
        8'b11111100,
        8'b00000100,
        8'b00000010,
        8'b11111101,
        8'b00000100,
        8'b11111110,
        8'b11111111,
        8'b00000010,
        8'b00000011,
        8'b00000101,
        8'b11111101,
        8'b00000001,
        8'b00000010,
        8'b00000001,
        8'b00000110,
        8'b00000100,
        8'b00000001,
        8'b00000101,
        8'b00000101,
        8'b00000110,
        8'b00000010,
        8'b11111010,
        8'b11111111,
        8'b11111100,
        8'b00000001,
        8'b11111100,
        8'b11110111,
        8'b00000010,
        8'b00000011,
        8'b00000101,
        8'b00001000,
        8'b11111101,
        8'b00000100,
        8'b00000010,
        8'b00000111,
        8'b11111101,
        8'b11111110,
        8'b11111010,
        8'b11111100,
        8'b00000110,
        8'b00000111,
        8'b00000001,
        8'b00001011,
        8'b00000001,
        8'b00000010,
        8'b11111001,
        8'b11111100,
        8'b11111100,
        8'b11111011,
        8'b11111110,
        8'b00000010,
        8'b11111111,
        8'b00000010,
        8'b11111111,
        8'b11111111,
        8'b00000101,
        8'b11111100,
        8'b00000111,
        8'b11111111,
        8'b11111010,
        8'b11111111,
        8'b00000001,
        8'b00000010,
        8'b00000100,
        8'b11111101,
        8'b00000100,
        8'b00000000,
        8'b00000101,
        8'b11111011,
        8'b11111010,
        8'b00000000,
        8'b00000001,
        8'b00000111,
        8'b00000010,
        8'b00000010,
        8'b00000001,
        8'b00000000,
        8'b11111011,
        8'b00000100,
        8'b11111100,
        8'b00000000,
        8'b11111111,
        8'b00000001,
        8'b11111100,
        8'b00000010,
        8'b11111100,
        8'b11111101,
        8'b00000100,
        8'b11111110,
        8'b11111101,
        8'b00000101,
        8'b00000100,
        8'b11111111,
        8'b11111010,
        8'b00000011,
        8'b11111101,
        8'b00000010,
        8'b11111011,
        8'b00000010,
        8'b00000001,
        8'b00000100,
        8'b00000010,
        8'b00000100,
        8'b11111111,
        8'b00000000,
        8'b11111111,
        8'b00000011,
        8'b00000000,
        8'b00000100,
        8'b00000000,
        8'b11111010,
        8'b00000011,
        8'b00000000,
        8'b11111111,
        8'b00000000,
        8'b00001000,
        8'b11111001,
        8'b00000001,
        8'b00000000,
        8'b11111111,
        8'b00001011,
        8'b00000100,
        8'b00000010,
        8'b00000001,
        8'b11111101,
        8'b00000100,
        8'b00000011,
        8'b11110110,
        8'b00000011,
        8'b11111011,
        8'b00000000,
        8'b00000110,
        8'b00000000,
        8'b00001000,
        8'b11111110,
        8'b11111111,
        8'b00000010,
        8'b00000011,
        8'b00000100,
        8'b11111011,
        8'b00000011,
        8'b00000101,
        8'b11111111,
        8'b00000000,
        8'b00000001,
        8'b11111111,
        8'b00000001,
        8'b00000010,
        8'b00000010,
        8'b11111100,
        8'b00000010,
        8'b00000100,
        8'b00000011,
        8'b00000011,
        8'b00000010,
        8'b00000000,
        8'b00000100,
        8'b00000000,
        8'b00000011,
        8'b00000100
    };
    assign values_bs = {
        8'b11111111,
        8'b11111100,
        8'b00000010,
        8'b11111110,
        8'b00000001,
        8'b11111100,
        8'b11111111,
        8'b00000010,
        8'b11111110,
        8'b11111110,
        8'b00000011,
        8'b00000001,
        8'b11111110,
        8'b00000100,
        8'b00000001,
        8'b11111110
    };
    assign values_wt = {
        8'b11111110,
        8'b11111110,
        8'b00000010,
        8'b00000101,
        8'b11111110,
        8'b00000110,
        8'b00000001,
        8'b11111101,
        8'b00000001,
        8'b11111010,
        8'b00000110,
        8'b00001101,
        8'b11111100,
        8'b11111100,
        8'b11110111,
        8'b11111001,
        8'b11111000,
        8'b00000001,
        8'b00000101,
        8'b00000111,
        8'b00001011,
        8'b11110010,
        8'b00001001,
        8'b00000001,
        8'b11111010,
        8'b11111111,
        8'b11111111,
        8'b11111101,
        8'b11111111,
        8'b11111010,
        8'b00000101,
        8'b11110001,
        8'b00000001,
        8'b11111100,
        8'b11111011,
        8'b11111010,
        8'b11110101,
        8'b11111101,
        8'b11111010,
        8'b00000011,
        8'b00000010,
        8'b11111000,
        8'b11111001,
        8'b11110100,
        8'b00000111,
        8'b11111011,
        8'b00001000,
        8'b00001101,
        8'b11111010,
        8'b00001000,
        8'b00001000,
        8'b00000101,
        8'b11111111,
        8'b11111100,
        8'b00000110,
        8'b11110111,
        8'b00000000,
        8'b11111010,
        8'b00000110,
        8'b00000100,
        8'b11111100,
        8'b11111110,
        8'b11111011,
        8'b11111010,
        8'b11111010,
        8'b00000101,
        8'b00000101,
        8'b00000000,
        8'b00000010,
        8'b00001000,
        8'b11111111,
        8'b11111111,
        8'b11111101,
        8'b00001100,
        8'b00000010,
        8'b00000100,
        8'b11111010,
        8'b00000001,
        8'b11111101,
        8'b00000100,
        8'b11111100,
        8'b11111001,
        8'b11111011,
        8'b11111010,
        8'b11111110,
        8'b11111011,
        8'b11111111,
        8'b00000011,
        8'b11111110,
        8'b11111010,
        8'b11111001,
        8'b00000000,
        8'b00000100,
        8'b11111101,
        8'b00000110,
        8'b11111011,
        8'b00000010,
        8'b11111100,
        8'b11111000,
        8'b11111001,
        8'b11110111,
        8'b00000111,
        8'b11111011,
        8'b00000011,
        8'b00000101,
        8'b00000100,
        8'b11110111,
        8'b00010000,
        8'b00001001,
        8'b00000010,
        8'b00001000,
        8'b00000110,
        8'b11111011,
        8'b11111110,
        8'b00000001,
        8'b11111101,
        8'b11111111,
        8'b00000000,
        8'b00000011,
        8'b11111101,
        8'b00000000,
        8'b00000110,
        8'b00000010,
        8'b00000010,
        8'b00000000,
        8'b11111101,
        8'b00000110,
        8'b00000001,
        8'b11111100,
        8'b00000011,
        8'b00000001,
        8'b11111111,
        8'b00000100,
        8'b11111101,
        8'b00000011,
        8'b11111100,
        8'b11111110,
        8'b11111100,
        8'b11111101,
        8'b11111001,
        8'b00000000,
        8'b11111100,
        8'b00000000,
        8'b11111111,
        8'b11111000,
        8'b00000001,
        8'b00000010,
        8'b11111101,
        8'b11111001,
        8'b00000001,
        8'b11111110,
        8'b11111011,
        8'b00000110,
        8'b00000001,
        8'b11111100,
        8'b00000010,
        8'b00000000,
        8'b11111100,
        8'b00001101,
        8'b11111111,
        8'b11111011,
        8'b11111101,
        8'b11111000,
        8'b11111100,
        8'b11111111,
        8'b00000011,
        8'b00000010,
        8'b00000101,
        8'b00000100,
        8'b00000101,
        8'b11111100,
        8'b11111000,
        8'b00000100,
        8'b00000111,
        8'b00000101,
        8'b00000010,
        8'b00000111,
        8'b11111100,
        8'b11110111,
        8'b11111111,
        8'b11111001,
        8'b00000010,
        8'b11111001,
        8'b00000111,
        8'b00001001,
        8'b11111010,
        8'b11110110,
        8'b00000000,
        8'b00001000,
        8'b00001000,
        8'b11110111,
        8'b00000110,
        8'b00000011,
        8'b00000110,
        8'b00001011,
        8'b00000010,
        8'b00000110,
        8'b00000110,
        8'b11111111,
        8'b11110101,
        8'b11110111,
        8'b11111110,
        8'b00000111,
        8'b00001000,
        8'b11110111,
        8'b11111100,
        8'b00000001,
        8'b00000100,
        8'b00000100,
        8'b11111101,
        8'b00000011,
        8'b11111111,
        8'b11111011,
        8'b11111110,
        8'b11111110,
        8'b11111101,
        8'b11111110,
        8'b00000001,
        8'b00000011,
        8'b00000000,
        8'b11111101,
        8'b00000001,
        8'b00000010,
        8'b11111110,
        8'b11111101,
        8'b00000001,
        8'b00000000,
        8'b00000010,
        8'b00000101,
        8'b11111101,
        8'b00000100,
        8'b11111100,
        8'b11110100,
        8'b00000001,
        8'b00000101,
        8'b11111110,
        8'b11111111,
        8'b11111101,
        8'b00000110,
        8'b00000000,
        8'b11111100,
        8'b00000100,
        8'b11111111,
        8'b00000101,
        8'b00000000,
        8'b00000001,
        8'b11111111,
        8'b00000010,
        8'b11111111,
        8'b00000100,
        8'b00000100,
        8'b00000001,
        8'b11111100,
        8'b00000000,
        8'b00000111,
        8'b00000001
    };
    assign mlp0_bs = {
        8'b11111110,
        8'b00000111,
        8'b00000001,
        8'b00000000,
        8'b00000100,
        8'b11111010,
        8'b11111111,
        8'b11111110,
        8'b00000100,
        8'b00000001,
        8'b11111111,
        8'b00000000,
        8'b00000010,
        8'b00000001,
        8'b00000010,
        8'b00000100
    };
    assign mlp0_wt = {
        8'b00000000,
        8'b11111010,
        8'b11111010,
        8'b00000000,
        8'b00000011,
        8'b00000000,
        8'b00001101,
        8'b00000001,
        8'b11111111,
        8'b00000101,
        8'b11111010,
        8'b11110100,
        8'b00000000,
        8'b00000011,
        8'b00000011,
        8'b00001000,
        8'b11111011,
        8'b00000100,
        8'b00000111,
        8'b00001101,
        8'b00000000,
        8'b11111100,
        8'b11111110,
        8'b11111101,
        8'b11111101,
        8'b11111011,
        8'b11111110,
        8'b00001100,
        8'b00000001,
        8'b00000000,
        8'b00000000,
        8'b00000010,
        8'b00000000,
        8'b11110100,
        8'b00000101,
        8'b00001100,
        8'b00000001,
        8'b11111100,
        8'b00010000,
        8'b00000001,
        8'b00000000,
        8'b11111111,
        8'b11111000,
        8'b00000100,
        8'b11111101,
        8'b00000011,
        8'b00000101,
        8'b00000010,
        8'b00000111,
        8'b11111000,
        8'b00000100,
        8'b00000111,
        8'b00000101,
        8'b00000110,
        8'b11111011,
        8'b00000100,
        8'b11111010,
        8'b00000100,
        8'b00000011,
        8'b11111011,
        8'b00000100,
        8'b11111000,
        8'b11111110,
        8'b00000011,
        8'b11110000,
        8'b00001010,
        8'b11111011,
        8'b00000101,
        8'b00000110,
        8'b11111111,
        8'b11111001,
        8'b11111011,
        8'b11111000,
        8'b11111110,
        8'b00000010,
        8'b00000000,
        8'b00000001,
        8'b11111100,
        8'b11111110,
        8'b00000011,
        8'b00000001,
        8'b11101110,
        8'b00001011,
        8'b00000111,
        8'b00001111,
        8'b11111010,
        8'b00001011,
        8'b00000011,
        8'b00000100,
        8'b00000110,
        8'b11110111,
        8'b11111101,
        8'b11111000,
        8'b00000110,
        8'b00000101,
        8'b11111101,
        8'b00000010,
        8'b11111110,
        8'b11111011,
        8'b11111111,
        8'b00000100,
        8'b00000101,
        8'b00001010,
        8'b00000101,
        8'b00000011,
        8'b00000100,
        8'b11110110,
        8'b00000011,
        8'b11111101,
        8'b00000100,
        8'b00000101,
        8'b00000111,
        8'b00000100,
        8'b00000100,
        8'b00000000,
        8'b00001001,
        8'b00000001,
        8'b00000110,
        8'b00001100,
        8'b11111111,
        8'b00000110,
        8'b00000101,
        8'b11111011,
        8'b11110001,
        8'b11111100,
        8'b00000101,
        8'b00000111,
        8'b11110100,
        8'b11111110,
        8'b00000010,
        8'b00000000,
        8'b00000100,
        8'b11111100,
        8'b11111100,
        8'b11111000,
        8'b00000001,
        8'b11111110,
        8'b00000100,
        8'b11111001,
        8'b00001100,
        8'b11111111,
        8'b11111110,
        8'b00000011,
        8'b00000001,
        8'b00000100,
        8'b11111011,
        8'b00000000,
        8'b00000110,
        8'b00000110,
        8'b11111011,
        8'b00000001,
        8'b00000011,
        8'b00000001,
        8'b00000100,
        8'b00000001,
        8'b00001010,
        8'b11111100,
        8'b00000001,
        8'b00000011,
        8'b00000001,
        8'b11111111,
        8'b11110101,
        8'b11110110,
        8'b11111010,
        8'b11110100,
        8'b11111110,
        8'b00000111,
        8'b00000101,
        8'b00000001,
        8'b11111011,
        8'b11111010,
        8'b00000001,
        8'b11111100,
        8'b00000011,
        8'b00000011,
        8'b11111110,
        8'b00000001,
        8'b11111101,
        8'b11111001,
        8'b11111101,
        8'b11110111,
        8'b11111110,
        8'b00000011,
        8'b00000001,
        8'b00000011,
        8'b11111101,
        8'b11111010,
        8'b00000101,
        8'b11111101,
        8'b00000010,
        8'b00000101,
        8'b00001001,
        8'b11111101,
        8'b00000111,
        8'b11111001,
        8'b00001010,
        8'b00000100,
        8'b00001010,
        8'b00000100,
        8'b11110000,
        8'b11111110,
        8'b00000001,
        8'b00000110,
        8'b00001000,
        8'b00000001,
        8'b11111111,
        8'b11111110,
        8'b00000000,
        8'b00000110,
        8'b00000001,
        8'b11111001,
        8'b11111110,
        8'b00001000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000011,
        8'b00001001,
        8'b11110111,
        8'b00001001,
        8'b11111100,
        8'b11111111,
        8'b00000101,
        8'b00000111,
        8'b11111100,
        8'b00000011,
        8'b11111010,
        8'b11111111,
        8'b00000000,
        8'b00000111,
        8'b11110011,
        8'b00000011,
        8'b11111010,
        8'b11110000,
        8'b00000001,
        8'b00001011,
        8'b00000000,
        8'b11111011,
        8'b11111011,
        8'b00000001,
        8'b11110111,
        8'b11111011,
        8'b00000001,
        8'b11110010,
        8'b00000110,
        8'b00001100,
        8'b11111111,
        8'b00000101,
        8'b00000001,
        8'b00000100,
        8'b11111110,
        8'b11111010,
        8'b11111110,
        8'b11111110,
        8'b00000001,
        8'b00000100
    };
    assign mlp1_bs = {
        8'b11111110,
        8'b11111111,
        8'b00000001,
        8'b11111111,
        8'b11111010,
        8'b00000001,
        8'b00000011,
        8'b00000010,
        8'b00000000,
        8'b11111111,
        8'b00000000,
        8'b11111111,
        8'b00000000,
        8'b11111111,
        8'b11111101,
        8'b11111111
    };
    assign mlp1_wt = {
        8'b00000001,
        8'b11111110,
        8'b00000011,
        8'b00000001,
        8'b11110111,
        8'b00000100,
        8'b00000010,
        8'b11111010,
        8'b00000010,
        8'b00001010,
        8'b11111100,
        8'b11111010,
        8'b00000111,
        8'b11111111,
        8'b00000010,
        8'b00000011,
        8'b11111111,
        8'b11111101,
        8'b11110111,
        8'b11111010,
        8'b00001101,
        8'b00000101,
        8'b00000011,
        8'b11111100,
        8'b11111111,
        8'b11111001,
        8'b00000011,
        8'b00000010,
        8'b00000001,
        8'b00000101,
        8'b11111111,
        8'b11111010,
        8'b00000111,
        8'b11111110,
        8'b11111100,
        8'b00000100,
        8'b11111001,
        8'b00000011,
        8'b00000010,
        8'b11111100,
        8'b11111110,
        8'b11111011,
        8'b11111011,
        8'b00000100,
        8'b11110110,
        8'b00000011,
        8'b00000101,
        8'b11111000,
        8'b11111011,
        8'b00000111,
        8'b00000011,
        8'b11111011,
        8'b00000001,
        8'b00000001,
        8'b11111101,
        8'b00001000,
        8'b00000000,
        8'b00000001,
        8'b11111101,
        8'b11111110,
        8'b00000001,
        8'b11111100,
        8'b00000101,
        8'b00000001,
        8'b00000111,
        8'b11110111,
        8'b00000000,
        8'b00000111,
        8'b11110110,
        8'b00000001,
        8'b00000011,
        8'b11111001,
        8'b11111111,
        8'b00000010,
        8'b11111100,
        8'b00000001,
        8'b11111010,
        8'b00000100,
        8'b00000011,
        8'b11111110,
        8'b00000001,
        8'b00000011,
        8'b11111100,
        8'b11111100,
        8'b00000010,
        8'b00000110,
        8'b11111110,
        8'b00000010,
        8'b11111110,
        8'b11111001,
        8'b11111100,
        8'b11111111,
        8'b11111101,
        8'b00000010,
        8'b00000101,
        8'b11111011,
        8'b11111110,
        8'b00000010,
        8'b00000011,
        8'b11111111,
        8'b00000011,
        8'b11111001,
        8'b00000000,
        8'b00000010,
        8'b00000101,
        8'b00000010,
        8'b00000110,
        8'b11111110,
        8'b00000001,
        8'b11111100,
        8'b11111010,
        8'b00000111,
        8'b00000110,
        8'b11111010,
        8'b00000001,
        8'b00001010,
        8'b11111101,
        8'b11111001,
        8'b00000111,
        8'b11110110,
        8'b11111100,
        8'b00000001,
        8'b00000101,
        8'b00000011,
        8'b11111001,
        8'b00000101,
        8'b11111010,
        8'b11111101,
        8'b00000100,
        8'b11111110,
        8'b00000010,
        8'b00000100,
        8'b11111111,
        8'b11110110,
        8'b00000110,
        8'b11111010,
        8'b11111110,
        8'b11111110,
        8'b00001001,
        8'b00000010,
        8'b11111001,
        8'b00000100,
        8'b11111010,
        8'b00000001,
        8'b00000101,
        8'b11111001,
        8'b00000000,
        8'b00000100,
        8'b00000010,
        8'b11111011,
        8'b00000001,
        8'b11111000,
        8'b00000010,
        8'b00000001,
        8'b00000101,
        8'b00000111,
        8'b11111111,
        8'b00000011,
        8'b11111001,
        8'b00000010,
        8'b11111100,
        8'b00000110,
        8'b00000000,
        8'b11111111,
        8'b11111111,
        8'b00000011,
        8'b11111111,
        8'b00000111,
        8'b11111110,
        8'b11111111,
        8'b11111011,
        8'b11111110,
        8'b11111101,
        8'b11111110,
        8'b00000111,
        8'b11111100,
        8'b11111111,
        8'b11111101,
        8'b11111111,
        8'b11111111,
        8'b11111010,
        8'b00000100,
        8'b00000010,
        8'b11111100,
        8'b00000011,
        8'b00000110,
        8'b11111110,
        8'b11111111,
        8'b00001101,
        8'b11111100,
        8'b00000001,
        8'b00000001,
        8'b11111111,
        8'b00000101,
        8'b11111101,
        8'b11111001,
        8'b00000010,
        8'b00001010,
        8'b11111001,
        8'b00000111,
        8'b00000100,
        8'b11111101,
        8'b11111011,
        8'b11111010,
        8'b00000111,
        8'b11111110,
        8'b00000100,
        8'b00000011,
        8'b00000011,
        8'b11111010,
        8'b00000100,
        8'b00001001,
        8'b11111100,
        8'b11111000,
        8'b00000010,
        8'b11111011,
        8'b00000001,
        8'b11111111,
        8'b00000101,
        8'b00000101,
        8'b11111010,
        8'b00000010,
        8'b11111000,
        8'b00000100,
        8'b00000011,
        8'b11110111,
        8'b11111011,
        8'b00000010,
        8'b11111011,
        8'b00000010,
        8'b00000110,
        8'b11110110,
        8'b00000000,
        8'b11111111,
        8'b11111111,
        8'b00000110,
        8'b00000101,
        8'b00000011,
        8'b11111101,
        8'b11111101,
        8'b00000000,
        8'b00000100,
        8'b00001000,
        8'b00000111,
        8'b11111011,
        8'b11111111,
        8'b00000011,
        8'b00000011,
        8'b00000001,
        8'b11111101,
        8'b11111010,
        8'b11111101,
        8'b11110001,
        8'b11111011,
        8'b00000011,
        8'b00000001
    };
    assign ps_wt = {
        8'b00001100,
        8'b00000000,
        8'b11101000,
        8'b11101110,
        8'b00000111,
        8'b11111001,
        8'b00001100,
        8'b00011100,
        8'b00011001,
        8'b11111111,
        8'b00001010,
        8'b00001010,
        8'b11100111,
        8'b00001000,
        8'b11101001,
        8'b11110001,
        8'b00010001,
        8'b11110111,
        8'b11111100,
        8'b00001100,
        8'b00000110,
        8'b11011011,
        8'b11111011,
        8'b11111011,
        8'b11110000,
        8'b11100100,
        8'b11111000,
        8'b00001000,
        8'b00001001,
        8'b00000100,
        8'b11110101,
        8'b00000001,
        8'b00000011,
        8'b11100001,
        8'b00101010,
        8'b11111001,
        8'b11101000,
        8'b11110000,
        8'b11011100,
        8'b00000101,
        8'b11111001,
        8'b11100101,
        8'b11110110,
        8'b11110011,
        8'b00001101,
        8'b00010111,
        8'b00100000,
        8'b11101010,
        8'b00001100,
        8'b00011101,
        8'b00010110,
        8'b00000100,
        8'b11111011,
        8'b00000101,
        8'b11101010,
        8'b00010000,
        8'b00000100,
        8'b00001100,
        8'b00100011,
        8'b00010000,
        8'b11110000,
        8'b00000000,
        8'b00000110,
        8'b00010110,
        8'b00001000,
        8'b11110010,
        8'b00000011,
        8'b00000100,
        8'b11100100,
        8'b00010010,
        8'b00001100,
        8'b00000001,
        8'b00000001,
        8'b00000001,
        8'b00001100,
        8'b00001101,
        8'b00010100,
        8'b00001010,
        8'b11100010,
        8'b11110111,
        8'b11100011,
        8'b00000000,
        8'b11111100,
        8'b11111111,
        8'b00010111,
        8'b11011000,
        8'b00100010,
        8'b00110100,
        8'b11111000,
        8'b00000101,
        8'b00000110,
        8'b11101011,
        8'b00001001,
        8'b00001001,
        8'b00010000,
        8'b11111110,
        8'b00000010,
        8'b00010100,
        8'b00011001,
        8'b00001110,
        8'b00010000,
        8'b11110111,
        8'b11010111,
        8'b00000101,
        8'b00010101,
        8'b00100001,
        8'b11101101,
        8'b00001101,
        8'b00001111,
        8'b11110110,
        8'b00000000,
        8'b00010111,
        8'b11110001,
        8'b11101110,
        8'b11110101,
        8'b00010110,
        8'b00000100,
        8'b11111001,
        8'b00000000,
        8'b11111101,
        8'b00011010,
        8'b00010100,
        8'b11111111,
        8'b00000000,
        8'b00000001,
        8'b00010000,
        8'b00011001,
        8'b11111000,
        8'b00010100,
        8'b11111010,
        8'b00001000,
        8'b11110010,
        8'b00001000,
        8'b11101111,
        8'b11111011,
        8'b11110001,
        8'b00110001,
        8'b00010101,
        8'b00001011,
        8'b00000001,
        8'b11111101,
        8'b00011000,
        8'b11011111,
        8'b00100000,
        8'b11111111,
        8'b11111101,
        8'b00000001,
        8'b00010100,
        8'b11111011,
        8'b11101100,
        8'b11011010,
        8'b11110100,
        8'b00000010,
        8'b00010011,
        8'b11100101,
        8'b11100011,
        8'b00000011,
        8'b11111100,
        8'b11111001,
        8'b00001000,
        8'b11011101,
        8'b11100100,
        8'b11110011,
        8'b11101111,
        8'b11111100,
        8'b11110001,
        8'b11110000,
        8'b00011000,
        8'b11110110,
        8'b11100110,
        8'b11100100,
        8'b00000011,
        8'b00011100,
        8'b11101111,
        8'b00000010,
        8'b00010101,
        8'b11111010,
        8'b00010001,
        8'b11110011,
        8'b11111111,
        8'b11011100,
        8'b00011011,
        8'b11111101,
        8'b00010011,
        8'b11111111,
        8'b00001101,
        8'b11110001,
        8'b11101110,
        8'b11111110,
        8'b00010100,
        8'b00000011,
        8'b11110101,
        8'b11110110,
        8'b00010111,
        8'b11101101,
        8'b11110111,
        8'b00000110,
        8'b00011000,
        8'b00010011,
        8'b11110000,
        8'b11110010,
        8'b11111010,
        8'b11101001,
        8'b00000111,
        8'b11101100,
        8'b00000001,
        8'b11111111,
        8'b00010001,
        8'b11110101,
        8'b11111101,
        8'b00100000,
        8'b11100010,
        8'b00001010,
        8'b11101111,
        8'b00010000,
        8'b11111111,
        8'b11101001,
        8'b00011001,
        8'b11101001,
        8'b00001100,
        8'b11110011,
        8'b00001001,
        8'b11110011,
        8'b00010011,
        8'b11110010,
        8'b11110001,
        8'b11110100,
        8'b00010010,
        8'b11100101,
        8'b00000100,
        8'b00010101,
        8'b11110010,
        8'b11111110,
        8'b00010011,
        8'b11110110,
        8'b11100111,
        8'b00001111,
        8'b00011111,
        8'b11101100,
        8'b11100111,
        8'b00100001,
        8'b00101111,
        8'b11011110,
        8'b00011001,
        8'b11111000,
        8'b00000011,
        8'b00010110,
        8'b00001000,
        8'b00001111,
        8'b00011000,
        8'b11111000,
        8'b11110100,
        8'b00011001,
        8'b11111011,
        8'b00011010,
        8'b00001011
    };


    // State machine
    typedef enum {
        IDLE,
        READ_CLASSIFIER_BS,
        READ_CLASSIFIER_WT,
        READ_EMBEDDING_BS,
        READ_EMBEDDING_WT,
        READ_CLS_TOKEN_WT,
        READ_FINAL_BS,
        READ_FINAL_WT,
        READ_KEYS_BS,
        READ_KEYS_WT,
        READ_QUERIES_BS,
        READ_QUERIES_WT,
        READ_VALUES_BS,
        READ_VALUES_WT,
        READ_MLP0_BS,
        READ_MLP0_WT,
        READ_MLP1_BS,
        READ_MLP1_WT,
        READ_PS_WT
    } state_t;
    state_t state, next_state;

    // State register
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
        end else begin
            state <= next_state;
        end
    end

    // Next state logic
    always_comb begin
        case (state)
            IDLE: begin
                if (start) begin
                    case (addr)
                        8'h01:   next_state = READ_CLASSIFIER_BS;
                        8'h02:   next_state = READ_CLASSIFIER_WT;
                        8'h03:   next_state = READ_EMBEDDING_BS;
                        8'h04:   next_state = READ_EMBEDDING_WT;
                        8'h05:   next_state = READ_CLS_TOKEN_WT;
                        8'h06:   next_state = READ_FINAL_BS;
                        8'h07:   next_state = READ_FINAL_WT;
                        8'h08:   next_state = READ_KEYS_BS;
                        8'h09:   next_state = READ_KEYS_WT;
                        8'h0A:   next_state = READ_QUERIES_BS;
                        8'h0B:   next_state = READ_QUERIES_WT;
                        8'h0C:   next_state = READ_VALUES_BS;
                        8'h0D:   next_state = READ_VALUES_WT;
                        8'h0E:   next_state = READ_MLP0_BS;
                        8'h0F:   next_state = READ_MLP0_WT;
                        8'h10:   next_state = READ_MLP1_BS;
                        8'h11:   next_state = READ_MLP1_WT;
                        8'h12:   next_state = READ_PS_WT;
                        default: next_state = IDLE;
                    endcase
                end else begin
                    next_state = state;
                end
            end
            READ_CLASSIFIER_BS: begin
                if (array_index == CLASSIFIER_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_CLASSIFIER_WT: begin
                if (array_index == CLASSIFIER_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_EMBEDDING_BS: begin
                if (array_index == EMBEDDING_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_EMBEDDING_WT: begin
                if (array_index == EMBEDDING_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_CLS_TOKEN_WT: begin
                if (array_index == CLS_TOKEN_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_FINAL_BS: begin
                if (array_index == FINAL_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_FINAL_WT: begin
                if (array_index == FINAL_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_KEYS_BS: begin
                if (array_index == KEYS_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_KEYS_WT: begin
                if (array_index == KEYS_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_QUERIES_BS: begin
                if (array_index == QUERIES_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_QUERIES_WT: begin
                if (array_index == QUERIES_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_VALUES_BS: begin
                if (array_index == VALUES_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_VALUES_WT: begin
                if (array_index == VALUES_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_MLP0_BS: begin
                if (array_index == MLP0_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_MLP0_WT: begin
                if (array_index == MLP0_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_MLP1_BS: begin
                if (array_index == MLP1_BS_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_MLP1_WT: begin
                if (array_index == MLP1_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            READ_PS_WT: begin
                if (array_index == PS_WT_CNT) begin
                    next_state = IDLE;
                end else begin
                    next_state = state;
                end
            end
            default: begin
                next_state = state;
            end
        endcase
    end


    // Array index logic
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            array_index <= '0;
        end else begin
            array_index <= array_index_ns;
        end
    end

    // array index 
    always_comb begin
        if (rst) begin
            array_index_ns = '0;
        end else begin
            case (state)
                IDLE: begin
                    array_index_ns = '0;
                end
                READ_CLASSIFIER_BS: begin
                    if (array_index == CLASSIFIER_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_CLASSIFIER_WT: begin
                    if (array_index == CLASSIFIER_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_EMBEDDING_BS: begin
                    if (array_index == EMBEDDING_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_EMBEDDING_WT: begin
                    if (array_index == EMBEDDING_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_CLS_TOKEN_WT: begin
                    if (array_index == CLS_TOKEN_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_FINAL_BS: begin
                    if (array_index == FINAL_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_FINAL_WT: begin
                    if (array_index == FINAL_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_KEYS_BS: begin
                    if (array_index == KEYS_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_KEYS_WT: begin
                    if (array_index == KEYS_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_QUERIES_BS: begin
                    if (array_index == QUERIES_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_QUERIES_WT: begin
                    if (array_index == QUERIES_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_VALUES_BS: begin
                    if (array_index == VALUES_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_VALUES_WT: begin
                    if (array_index == VALUES_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_MLP0_BS: begin
                    if (array_index == MLP0_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_MLP0_WT: begin
                    if (array_index == MLP0_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_MLP1_BS: begin
                    if (array_index == MLP1_BS_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_MLP1_WT: begin
                    if (array_index == MLP1_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                READ_PS_WT: begin
                    if (array_index == PS_WT_CNT) begin
                        array_index_ns = 0;
                    end else begin
                        array_index_ns = array_index + 1;
                    end
                end
                default: begin
                    array_index_ns = array_index + 1;
                end
            endcase
        end
    end


    // done logic 
    always_comb begin
        done = 1'b0;
        case (state)
            READ_CLASSIFIER_BS: begin
                data = classifier_bs[array_index];
                if (array_index == 6) begin
                    done = 1'b1;
                end
            end
            READ_CLASSIFIER_WT: begin
                data = classifier_wt[array_index];
                if (array_index == 96) begin
                    done = 1'b1;
                end
            end
            READ_EMBEDDING_BS: begin
                data = embedding_bs[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_EMBEDDING_WT: begin
                data = embedding_wt[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_CLS_TOKEN_WT: begin
                data = cls_token_wt[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_FINAL_BS: begin
                data = final_bs[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_FINAL_WT: begin
                data = final_wt[array_index];
                if (array_index == 256) begin
                    done = 1'b1;
                end
            end
            READ_KEYS_BS: begin
                data = keys_bs[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_KEYS_WT: begin
                data = keys_wt[array_index];
                if (array_index == 256) begin
                    done = 1'b1;
                end
            end
            READ_QUERIES_BS: begin
                data = queries_bs[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_QUERIES_WT: begin
                data = queries_wt[array_index];
                if (array_index == 256) begin
                    done = 1'b1;
                end
            end
            READ_VALUES_BS: begin
                data = values_bs[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_VALUES_WT: begin
                data = values_wt[array_index];
                if (array_index == 256) begin
                    done = 1'b1;
                end
            end
            READ_MLP0_BS: begin
                data = mlp0_bs[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_MLP0_WT: begin
                data = mlp0_wt[array_index];
                if (array_index == 256) begin
                    done = 1'b1;
                end
            end
            READ_MLP1_BS: begin
                data = mlp1_bs[array_index];
                if (array_index == 16) begin
                    done = 1'b1;
                end
            end
            READ_MLP1_WT: begin
                data = mlp1_wt[array_index];
                if (array_index == 256) begin
                    done = 1'b1;
                end
            end
            READ_PS_WT: begin
                data = ps_wt[array_index];
                if (array_index == 256) begin
                    done = 1'b1;
                end
            end
            default: begin
                data = '0;
            end
        endcase
    end

    always_ff @(posedge clk, posedge rst) begin
        if (rst) data_o <= 0;
        else if (next_state == IDLE) data_o <= data_o;
        else data_o <= data;
    end

endmodule
